show_info_rom[542] = '{ v_ada: 10'd0, v_din_t: 0, adb_diff: 8'h00, vram_write: 0, mem_read: 1};
show_info_rom[544] = '{ v_ada: 10'd544, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[545] = '{ v_ada: 10'd545, v_din_t: 1, adb_diff: 8'h01, vram_write: 1, mem_read: 1};
show_info_rom[546] = '{ v_ada: 10'd546, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[547] = '{ v_ada: 10'd547, v_din_t: 1, adb_diff: 8'h02, vram_write: 1, mem_read: 1};
show_info_rom[548] = '{ v_ada: 10'd548, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[549] = '{ v_ada: 10'd549, v_din_t: 1, adb_diff: 8'h03, vram_write: 1, mem_read: 1};
show_info_rom[550] = '{ v_ada: 10'd550, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[551] = '{ v_ada: 10'd551, v_din_t: 1, adb_diff: 8'h04, vram_write: 1, mem_read: 1};
show_info_rom[553] = '{ v_ada: 10'd553, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[554] = '{ v_ada: 10'd554, v_din_t: 1, adb_diff: 8'h05, vram_write: 1, mem_read: 1};
show_info_rom[555] = '{ v_ada: 10'd555, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[556] = '{ v_ada: 10'd556, v_din_t: 1, adb_diff: 8'h06, vram_write: 1, mem_read: 1};
show_info_rom[557] = '{ v_ada: 10'd557, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[558] = '{ v_ada: 10'd558, v_din_t: 1, adb_diff: 8'h07, vram_write: 1, mem_read: 1};
show_info_rom[559] = '{ v_ada: 10'd559, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[560] = '{ v_ada: 10'd560, v_din_t: 1, adb_diff: 8'h08, vram_write: 1, mem_read: 1};
show_info_rom[563] = '{ v_ada: 10'd563, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[564] = '{ v_ada: 10'd564, v_din_t: 1, adb_diff: 8'h09, vram_write: 1, mem_read: 1};
show_info_rom[565] = '{ v_ada: 10'd565, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[566] = '{ v_ada: 10'd566, v_din_t: 1, adb_diff: 8'h0A, vram_write: 1, mem_read: 1};
show_info_rom[567] = '{ v_ada: 10'd567, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[568] = '{ v_ada: 10'd568, v_din_t: 1, adb_diff: 8'h0B, vram_write: 1, mem_read: 1};
show_info_rom[569] = '{ v_ada: 10'd569, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[570] = '{ v_ada: 10'd570, v_din_t: 1, adb_diff: 8'h0C, vram_write: 1, mem_read: 1};
show_info_rom[572] = '{ v_ada: 10'd572, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[573] = '{ v_ada: 10'd573, v_din_t: 1, adb_diff: 8'h0D, vram_write: 1, mem_read: 1};
show_info_rom[574] = '{ v_ada: 10'd574, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[575] = '{ v_ada: 10'd575, v_din_t: 1, adb_diff: 8'h0E, vram_write: 1, mem_read: 1};
show_info_rom[576] = '{ v_ada: 10'd576, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[577] = '{ v_ada: 10'd577, v_din_t: 1, adb_diff: 8'h0F, vram_write: 1, mem_read: 1};
show_info_rom[578] = '{ v_ada: 10'd578, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[579] = '{ v_ada: 10'd579, v_din_t: 1, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[602] = '{ v_ada: 10'd0, v_din_t: 0, adb_diff: 8'h10, vram_write: 0, mem_read: 1};
show_info_rom[604] = '{ v_ada: 10'd604, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[605] = '{ v_ada: 10'd605, v_din_t: 1, adb_diff: 8'h11, vram_write: 1, mem_read: 1};
show_info_rom[606] = '{ v_ada: 10'd606, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[607] = '{ v_ada: 10'd607, v_din_t: 1, adb_diff: 8'h12, vram_write: 1, mem_read: 1};
show_info_rom[608] = '{ v_ada: 10'd608, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[609] = '{ v_ada: 10'd609, v_din_t: 1, adb_diff: 8'h13, vram_write: 1, mem_read: 1};
show_info_rom[610] = '{ v_ada: 10'd610, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[611] = '{ v_ada: 10'd611, v_din_t: 1, adb_diff: 8'h14, vram_write: 1, mem_read: 1};
show_info_rom[613] = '{ v_ada: 10'd613, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[614] = '{ v_ada: 10'd614, v_din_t: 1, adb_diff: 8'h15, vram_write: 1, mem_read: 1};
show_info_rom[615] = '{ v_ada: 10'd615, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[616] = '{ v_ada: 10'd616, v_din_t: 1, adb_diff: 8'h16, vram_write: 1, mem_read: 1};
show_info_rom[617] = '{ v_ada: 10'd617, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[618] = '{ v_ada: 10'd618, v_din_t: 1, adb_diff: 8'h17, vram_write: 1, mem_read: 1};
show_info_rom[619] = '{ v_ada: 10'd619, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[620] = '{ v_ada: 10'd620, v_din_t: 1, adb_diff: 8'h18, vram_write: 1, mem_read: 1};
show_info_rom[623] = '{ v_ada: 10'd623, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[624] = '{ v_ada: 10'd624, v_din_t: 1, adb_diff: 8'h19, vram_write: 1, mem_read: 1};
show_info_rom[625] = '{ v_ada: 10'd625, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[626] = '{ v_ada: 10'd626, v_din_t: 1, adb_diff: 8'h1A, vram_write: 1, mem_read: 1};
show_info_rom[627] = '{ v_ada: 10'd627, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[628] = '{ v_ada: 10'd628, v_din_t: 1, adb_diff: 8'h1B, vram_write: 1, mem_read: 1};
show_info_rom[629] = '{ v_ada: 10'd629, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[630] = '{ v_ada: 10'd630, v_din_t: 1, adb_diff: 8'h1C, vram_write: 1, mem_read: 1};
show_info_rom[632] = '{ v_ada: 10'd632, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[633] = '{ v_ada: 10'd633, v_din_t: 1, adb_diff: 8'h1D, vram_write: 1, mem_read: 1};
show_info_rom[634] = '{ v_ada: 10'd634, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[635] = '{ v_ada: 10'd635, v_din_t: 1, adb_diff: 8'h1E, vram_write: 1, mem_read: 1};
show_info_rom[636] = '{ v_ada: 10'd636, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[637] = '{ v_ada: 10'd637, v_din_t: 1, adb_diff: 8'h1F, vram_write: 1, mem_read: 1};
show_info_rom[638] = '{ v_ada: 10'd638, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[639] = '{ v_ada: 10'd639, v_din_t: 1, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[662] = '{ v_ada: 10'd0, v_din_t: 0, adb_diff: 8'h20, vram_write: 0, mem_read: 1};
show_info_rom[664] = '{ v_ada: 10'd664, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[665] = '{ v_ada: 10'd665, v_din_t: 1, adb_diff: 8'h21, vram_write: 1, mem_read: 1};
show_info_rom[666] = '{ v_ada: 10'd666, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[667] = '{ v_ada: 10'd667, v_din_t: 1, adb_diff: 8'h22, vram_write: 1, mem_read: 1};
show_info_rom[668] = '{ v_ada: 10'd668, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[669] = '{ v_ada: 10'd669, v_din_t: 1, adb_diff: 8'h23, vram_write: 1, mem_read: 1};
show_info_rom[670] = '{ v_ada: 10'd670, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[671] = '{ v_ada: 10'd671, v_din_t: 1, adb_diff: 8'h24, vram_write: 1, mem_read: 1};
show_info_rom[673] = '{ v_ada: 10'd673, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[674] = '{ v_ada: 10'd674, v_din_t: 1, adb_diff: 8'h25, vram_write: 1, mem_read: 1};
show_info_rom[675] = '{ v_ada: 10'd675, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[676] = '{ v_ada: 10'd676, v_din_t: 1, adb_diff: 8'h26, vram_write: 1, mem_read: 1};
show_info_rom[677] = '{ v_ada: 10'd677, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[678] = '{ v_ada: 10'd678, v_din_t: 1, adb_diff: 8'h27, vram_write: 1, mem_read: 1};
show_info_rom[679] = '{ v_ada: 10'd679, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[680] = '{ v_ada: 10'd680, v_din_t: 1, adb_diff: 8'h28, vram_write: 1, mem_read: 1};
show_info_rom[683] = '{ v_ada: 10'd683, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[684] = '{ v_ada: 10'd684, v_din_t: 1, adb_diff: 8'h29, vram_write: 1, mem_read: 1};
show_info_rom[685] = '{ v_ada: 10'd685, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[686] = '{ v_ada: 10'd686, v_din_t: 1, adb_diff: 8'h2A, vram_write: 1, mem_read: 1};
show_info_rom[687] = '{ v_ada: 10'd687, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[688] = '{ v_ada: 10'd688, v_din_t: 1, adb_diff: 8'h2B, vram_write: 1, mem_read: 1};
show_info_rom[689] = '{ v_ada: 10'd689, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[690] = '{ v_ada: 10'd690, v_din_t: 1, adb_diff: 8'h2C, vram_write: 1, mem_read: 1};
show_info_rom[692] = '{ v_ada: 10'd692, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[693] = '{ v_ada: 10'd693, v_din_t: 1, adb_diff: 8'h2D, vram_write: 1, mem_read: 1};
show_info_rom[694] = '{ v_ada: 10'd694, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[695] = '{ v_ada: 10'd695, v_din_t: 1, adb_diff: 8'h2E, vram_write: 1, mem_read: 1};
show_info_rom[696] = '{ v_ada: 10'd696, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[697] = '{ v_ada: 10'd697, v_din_t: 1, adb_diff: 8'h2F, vram_write: 1, mem_read: 1};
show_info_rom[698] = '{ v_ada: 10'd698, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[699] = '{ v_ada: 10'd699, v_din_t: 1, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[722] = '{ v_ada: 10'd0, v_din_t: 0, adb_diff: 8'h30, vram_write: 0, mem_read: 1};
show_info_rom[724] = '{ v_ada: 10'd724, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[725] = '{ v_ada: 10'd725, v_din_t: 1, adb_diff: 8'h31, vram_write: 1, mem_read: 1};
show_info_rom[726] = '{ v_ada: 10'd726, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[727] = '{ v_ada: 10'd727, v_din_t: 1, adb_diff: 8'h32, vram_write: 1, mem_read: 1};
show_info_rom[728] = '{ v_ada: 10'd728, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[729] = '{ v_ada: 10'd729, v_din_t: 1, adb_diff: 8'h33, vram_write: 1, mem_read: 1};
show_info_rom[730] = '{ v_ada: 10'd730, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[731] = '{ v_ada: 10'd731, v_din_t: 1, adb_diff: 8'h34, vram_write: 1, mem_read: 1};
show_info_rom[733] = '{ v_ada: 10'd733, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[734] = '{ v_ada: 10'd734, v_din_t: 1, adb_diff: 8'h35, vram_write: 1, mem_read: 1};
show_info_rom[735] = '{ v_ada: 10'd735, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[736] = '{ v_ada: 10'd736, v_din_t: 1, adb_diff: 8'h36, vram_write: 1, mem_read: 1};
show_info_rom[737] = '{ v_ada: 10'd737, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[738] = '{ v_ada: 10'd738, v_din_t: 1, adb_diff: 8'h37, vram_write: 1, mem_read: 1};
show_info_rom[739] = '{ v_ada: 10'd739, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[740] = '{ v_ada: 10'd740, v_din_t: 1, adb_diff: 8'h38, vram_write: 1, mem_read: 1};
show_info_rom[743] = '{ v_ada: 10'd743, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[744] = '{ v_ada: 10'd744, v_din_t: 1, adb_diff: 8'h39, vram_write: 1, mem_read: 1};
show_info_rom[745] = '{ v_ada: 10'd745, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[746] = '{ v_ada: 10'd746, v_din_t: 1, adb_diff: 8'h3A, vram_write: 1, mem_read: 1};
show_info_rom[747] = '{ v_ada: 10'd747, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[748] = '{ v_ada: 10'd748, v_din_t: 1, adb_diff: 8'h3B, vram_write: 1, mem_read: 1};
show_info_rom[749] = '{ v_ada: 10'd749, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[750] = '{ v_ada: 10'd750, v_din_t: 1, adb_diff: 8'h3C, vram_write: 1, mem_read: 1};
show_info_rom[752] = '{ v_ada: 10'd752, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[753] = '{ v_ada: 10'd753, v_din_t: 1, adb_diff: 8'h3D, vram_write: 1, mem_read: 1};
show_info_rom[754] = '{ v_ada: 10'd754, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[755] = '{ v_ada: 10'd755, v_din_t: 1, adb_diff: 8'h3E, vram_write: 1, mem_read: 1};
show_info_rom[756] = '{ v_ada: 10'd756, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[757] = '{ v_ada: 10'd757, v_din_t: 1, adb_diff: 8'h3F, vram_write: 1, mem_read: 1};
show_info_rom[758] = '{ v_ada: 10'd758, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[759] = '{ v_ada: 10'd759, v_din_t: 1, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[782] = '{ v_ada: 10'd0, v_din_t: 0, adb_diff: 8'h40, vram_write: 0, mem_read: 1};
show_info_rom[784] = '{ v_ada: 10'd784, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[785] = '{ v_ada: 10'd785, v_din_t: 1, adb_diff: 8'h41, vram_write: 1, mem_read: 1};
show_info_rom[786] = '{ v_ada: 10'd786, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[787] = '{ v_ada: 10'd787, v_din_t: 1, adb_diff: 8'h42, vram_write: 1, mem_read: 1};
show_info_rom[788] = '{ v_ada: 10'd788, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[789] = '{ v_ada: 10'd789, v_din_t: 1, adb_diff: 8'h43, vram_write: 1, mem_read: 1};
show_info_rom[790] = '{ v_ada: 10'd790, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[791] = '{ v_ada: 10'd791, v_din_t: 1, adb_diff: 8'h44, vram_write: 1, mem_read: 1};
show_info_rom[793] = '{ v_ada: 10'd793, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[794] = '{ v_ada: 10'd794, v_din_t: 1, adb_diff: 8'h45, vram_write: 1, mem_read: 1};
show_info_rom[795] = '{ v_ada: 10'd795, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[796] = '{ v_ada: 10'd796, v_din_t: 1, adb_diff: 8'h46, vram_write: 1, mem_read: 1};
show_info_rom[797] = '{ v_ada: 10'd797, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[798] = '{ v_ada: 10'd798, v_din_t: 1, adb_diff: 8'h47, vram_write: 1, mem_read: 1};
show_info_rom[799] = '{ v_ada: 10'd799, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[800] = '{ v_ada: 10'd800, v_din_t: 1, adb_diff: 8'h48, vram_write: 1, mem_read: 1};
show_info_rom[803] = '{ v_ada: 10'd803, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[804] = '{ v_ada: 10'd804, v_din_t: 1, adb_diff: 8'h49, vram_write: 1, mem_read: 1};
show_info_rom[805] = '{ v_ada: 10'd805, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[806] = '{ v_ada: 10'd806, v_din_t: 1, adb_diff: 8'h4A, vram_write: 1, mem_read: 1};
show_info_rom[807] = '{ v_ada: 10'd807, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[808] = '{ v_ada: 10'd808, v_din_t: 1, adb_diff: 8'h4B, vram_write: 1, mem_read: 1};
show_info_rom[809] = '{ v_ada: 10'd809, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[810] = '{ v_ada: 10'd810, v_din_t: 1, adb_diff: 8'h4C, vram_write: 1, mem_read: 1};
show_info_rom[812] = '{ v_ada: 10'd812, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[813] = '{ v_ada: 10'd813, v_din_t: 1, adb_diff: 8'h4D, vram_write: 1, mem_read: 1};
show_info_rom[814] = '{ v_ada: 10'd814, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[815] = '{ v_ada: 10'd815, v_din_t: 1, adb_diff: 8'h4E, vram_write: 1, mem_read: 1};
show_info_rom[816] = '{ v_ada: 10'd816, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[817] = '{ v_ada: 10'd817, v_din_t: 1, adb_diff: 8'h4F, vram_write: 1, mem_read: 1};
show_info_rom[818] = '{ v_ada: 10'd818, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[819] = '{ v_ada: 10'd819, v_din_t: 1, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[842] = '{ v_ada: 10'd0, v_din_t: 0, adb_diff: 8'h50, vram_write: 0, mem_read: 1};
show_info_rom[844] = '{ v_ada: 10'd844, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[845] = '{ v_ada: 10'd845, v_din_t: 1, adb_diff: 8'h51, vram_write: 1, mem_read: 1};
show_info_rom[846] = '{ v_ada: 10'd846, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[847] = '{ v_ada: 10'd847, v_din_t: 1, adb_diff: 8'h52, vram_write: 1, mem_read: 1};
show_info_rom[848] = '{ v_ada: 10'd848, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[849] = '{ v_ada: 10'd849, v_din_t: 1, adb_diff: 8'h53, vram_write: 1, mem_read: 1};
show_info_rom[850] = '{ v_ada: 10'd850, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[851] = '{ v_ada: 10'd851, v_din_t: 1, adb_diff: 8'h54, vram_write: 1, mem_read: 1};
show_info_rom[853] = '{ v_ada: 10'd853, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[854] = '{ v_ada: 10'd854, v_din_t: 1, adb_diff: 8'h55, vram_write: 1, mem_read: 1};
show_info_rom[855] = '{ v_ada: 10'd855, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[856] = '{ v_ada: 10'd856, v_din_t: 1, adb_diff: 8'h56, vram_write: 1, mem_read: 1};
show_info_rom[857] = '{ v_ada: 10'd857, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[858] = '{ v_ada: 10'd858, v_din_t: 1, adb_diff: 8'h57, vram_write: 1, mem_read: 1};
show_info_rom[859] = '{ v_ada: 10'd859, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[860] = '{ v_ada: 10'd860, v_din_t: 1, adb_diff: 8'h58, vram_write: 1, mem_read: 1};
show_info_rom[863] = '{ v_ada: 10'd863, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[864] = '{ v_ada: 10'd864, v_din_t: 1, adb_diff: 8'h59, vram_write: 1, mem_read: 1};
show_info_rom[865] = '{ v_ada: 10'd865, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[866] = '{ v_ada: 10'd866, v_din_t: 1, adb_diff: 8'h5A, vram_write: 1, mem_read: 1};
show_info_rom[867] = '{ v_ada: 10'd867, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[868] = '{ v_ada: 10'd868, v_din_t: 1, adb_diff: 8'h5B, vram_write: 1, mem_read: 1};
show_info_rom[869] = '{ v_ada: 10'd869, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[870] = '{ v_ada: 10'd870, v_din_t: 1, adb_diff: 8'h5C, vram_write: 1, mem_read: 1};
show_info_rom[872] = '{ v_ada: 10'd872, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[873] = '{ v_ada: 10'd873, v_din_t: 1, adb_diff: 8'h5D, vram_write: 1, mem_read: 1};
show_info_rom[874] = '{ v_ada: 10'd874, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[875] = '{ v_ada: 10'd875, v_din_t: 1, adb_diff: 8'h5E, vram_write: 1, mem_read: 1};
show_info_rom[876] = '{ v_ada: 10'd876, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[877] = '{ v_ada: 10'd877, v_din_t: 1, adb_diff: 8'h5F, vram_write: 1, mem_read: 1};
show_info_rom[878] = '{ v_ada: 10'd878, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[879] = '{ v_ada: 10'd879, v_din_t: 1, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[902] = '{ v_ada: 10'd0, v_din_t: 0, adb_diff: 8'h60, vram_write: 0, mem_read: 1};
show_info_rom[904] = '{ v_ada: 10'd904, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[905] = '{ v_ada: 10'd905, v_din_t: 1, adb_diff: 8'h61, vram_write: 1, mem_read: 1};
show_info_rom[906] = '{ v_ada: 10'd906, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[907] = '{ v_ada: 10'd907, v_din_t: 1, adb_diff: 8'h62, vram_write: 1, mem_read: 1};
show_info_rom[908] = '{ v_ada: 10'd908, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[909] = '{ v_ada: 10'd909, v_din_t: 1, adb_diff: 8'h63, vram_write: 1, mem_read: 1};
show_info_rom[910] = '{ v_ada: 10'd910, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[911] = '{ v_ada: 10'd911, v_din_t: 1, adb_diff: 8'h64, vram_write: 1, mem_read: 1};
show_info_rom[913] = '{ v_ada: 10'd913, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[914] = '{ v_ada: 10'd914, v_din_t: 1, adb_diff: 8'h65, vram_write: 1, mem_read: 1};
show_info_rom[915] = '{ v_ada: 10'd915, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[916] = '{ v_ada: 10'd916, v_din_t: 1, adb_diff: 8'h66, vram_write: 1, mem_read: 1};
show_info_rom[917] = '{ v_ada: 10'd917, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[918] = '{ v_ada: 10'd918, v_din_t: 1, adb_diff: 8'h67, vram_write: 1, mem_read: 1};
show_info_rom[919] = '{ v_ada: 10'd919, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[920] = '{ v_ada: 10'd920, v_din_t: 1, adb_diff: 8'h68, vram_write: 1, mem_read: 1};
show_info_rom[923] = '{ v_ada: 10'd923, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[924] = '{ v_ada: 10'd924, v_din_t: 1, adb_diff: 8'h69, vram_write: 1, mem_read: 1};
show_info_rom[925] = '{ v_ada: 10'd925, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[926] = '{ v_ada: 10'd926, v_din_t: 1, adb_diff: 8'h6A, vram_write: 1, mem_read: 1};
show_info_rom[927] = '{ v_ada: 10'd927, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[928] = '{ v_ada: 10'd928, v_din_t: 1, adb_diff: 8'h6B, vram_write: 1, mem_read: 1};
show_info_rom[929] = '{ v_ada: 10'd929, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[930] = '{ v_ada: 10'd930, v_din_t: 1, adb_diff: 8'h6C, vram_write: 1, mem_read: 1};
show_info_rom[932] = '{ v_ada: 10'd932, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[933] = '{ v_ada: 10'd933, v_din_t: 1, adb_diff: 8'h6D, vram_write: 1, mem_read: 1};
show_info_rom[934] = '{ v_ada: 10'd934, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[935] = '{ v_ada: 10'd935, v_din_t: 1, adb_diff: 8'h6E, vram_write: 1, mem_read: 1};
show_info_rom[936] = '{ v_ada: 10'd936, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[937] = '{ v_ada: 10'd937, v_din_t: 1, adb_diff: 8'h6F, vram_write: 1, mem_read: 1};
show_info_rom[938] = '{ v_ada: 10'd938, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[939] = '{ v_ada: 10'd939, v_din_t: 1, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[962] = '{ v_ada: 10'd0, v_din_t: 0, adb_diff: 8'h70, vram_write: 0, mem_read: 1};
show_info_rom[964] = '{ v_ada: 10'd964, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[965] = '{ v_ada: 10'd965, v_din_t: 1, adb_diff: 8'h71, vram_write: 1, mem_read: 1};
show_info_rom[966] = '{ v_ada: 10'd966, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[967] = '{ v_ada: 10'd967, v_din_t: 1, adb_diff: 8'h72, vram_write: 1, mem_read: 1};
show_info_rom[968] = '{ v_ada: 10'd968, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[969] = '{ v_ada: 10'd969, v_din_t: 1, adb_diff: 8'h73, vram_write: 1, mem_read: 1};
show_info_rom[970] = '{ v_ada: 10'd970, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[971] = '{ v_ada: 10'd971, v_din_t: 1, adb_diff: 8'h74, vram_write: 1, mem_read: 1};
show_info_rom[973] = '{ v_ada: 10'd973, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[974] = '{ v_ada: 10'd974, v_din_t: 1, adb_diff: 8'h75, vram_write: 1, mem_read: 1};
show_info_rom[975] = '{ v_ada: 10'd975, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[976] = '{ v_ada: 10'd976, v_din_t: 1, adb_diff: 8'h76, vram_write: 1, mem_read: 1};
show_info_rom[977] = '{ v_ada: 10'd977, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[978] = '{ v_ada: 10'd978, v_din_t: 1, adb_diff: 8'h77, vram_write: 1, mem_read: 1};
show_info_rom[979] = '{ v_ada: 10'd979, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[980] = '{ v_ada: 10'd980, v_din_t: 1, adb_diff: 8'h78, vram_write: 1, mem_read: 1};
show_info_rom[983] = '{ v_ada: 10'd983, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[984] = '{ v_ada: 10'd984, v_din_t: 1, adb_diff: 8'h79, vram_write: 1, mem_read: 1};
show_info_rom[985] = '{ v_ada: 10'd985, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[986] = '{ v_ada: 10'd986, v_din_t: 1, adb_diff: 8'h7A, vram_write: 1, mem_read: 1};
show_info_rom[987] = '{ v_ada: 10'd987, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[988] = '{ v_ada: 10'd988, v_din_t: 1, adb_diff: 8'h7B, vram_write: 1, mem_read: 1};
show_info_rom[989] = '{ v_ada: 10'd989, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[990] = '{ v_ada: 10'd990, v_din_t: 1, adb_diff: 8'h7C, vram_write: 1, mem_read: 1};
show_info_rom[992] = '{ v_ada: 10'd992, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[993] = '{ v_ada: 10'd993, v_din_t: 1, adb_diff: 8'h7D, vram_write: 1, mem_read: 1};
show_info_rom[994] = '{ v_ada: 10'd994, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[995] = '{ v_ada: 10'd995, v_din_t: 1, adb_diff: 8'h7E, vram_write: 1, mem_read: 1};
show_info_rom[996] = '{ v_ada: 10'd996, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[997] = '{ v_ada: 10'd997, v_din_t: 1, adb_diff: 8'h7F, vram_write: 1, mem_read: 1};
show_info_rom[998] = '{ v_ada: 10'd998, v_din_t: 0, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[999] = '{ v_ada: 10'd999, v_din_t: 1, adb_diff: 8'h00, vram_write: 1, mem_read: 0};
