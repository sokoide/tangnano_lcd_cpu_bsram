902: begin adb <= operands[15:0] + 8'h60 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
904: begin v_ada <= 904; v_din <= to_hexchar(dout[7:4]); end
905: begin v_ada <= 905; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h61 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
906: begin v_ada <= 906; v_din <= to_hexchar(dout[7:4]); end
907: begin v_ada <= 907; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h62 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
908: begin v_ada <= 908; v_din <= to_hexchar(dout[7:4]); end
909: begin v_ada <= 909; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h63 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
910: begin v_ada <= 910; v_din <= to_hexchar(dout[7:4]); end
911: begin v_ada <= 911; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h64 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
913: begin v_ada <= 913; v_din <= to_hexchar(dout[7:4]); end
914: begin v_ada <= 914; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h65 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
915: begin v_ada <= 915; v_din <= to_hexchar(dout[7:4]); end
916: begin v_ada <= 916; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h66 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
917: begin v_ada <= 917; v_din <= to_hexchar(dout[7:4]); end
918: begin v_ada <= 918; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h67 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
919: begin v_ada <= 919; v_din <= to_hexchar(dout[7:4]); end
920: begin v_ada <= 920; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h68 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
923: begin v_ada <= 923; v_din <= to_hexchar(dout[7:4]); end
924: begin v_ada <= 924; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h69 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
925: begin v_ada <= 925; v_din <= to_hexchar(dout[7:4]); end
926: begin v_ada <= 926; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h6A & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
927: begin v_ada <= 927; v_din <= to_hexchar(dout[7:4]); end
928: begin v_ada <= 928; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h6B & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
929: begin v_ada <= 929; v_din <= to_hexchar(dout[7:4]); end
930: begin v_ada <= 930; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h6C & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
932: begin v_ada <= 932; v_din <= to_hexchar(dout[7:4]); end
933: begin v_ada <= 933; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h6D & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
934: begin v_ada <= 934; v_din <= to_hexchar(dout[7:4]); end
935: begin v_ada <= 935; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h6E & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
936: begin v_ada <= 936; v_din <= to_hexchar(dout[7:4]); end
937: begin v_ada <= 937; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h6F & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
938: begin v_ada <= 938; v_din <= to_hexchar(dout[7:4]); end
939: begin v_ada <= 939; v_din <= to_hexchar(dout[3:0]); end
