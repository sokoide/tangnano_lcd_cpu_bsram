//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Mon Apr  7 00:05:13 2025

module Gowin_pROM_font (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h000088C888C88000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h000000000000000000002C4C228880000004AA40084200000000088880088000;
defparam prom_inst_0.INIT_RAM_0A = 256'h000000008000000000000080C080000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000008800000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h00008444484448000000C00000844800000000000000000000008444444C4800;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000008444C0000008444480008000000844448000C0000008888C8888800;
defparam prom_inst_0.INIT_RAM_0E = 256'h00000000000000000000000000000000000084444C4448000000844448444800;
defparam prom_inst_0.INIT_RAM_0F = 256'h000000000844480000000000800000000000000C0C0000000000800000008000;
defparam prom_inst_0.INIT_RAM_10 = 256'h0000840000004800000084444844480000004444C44448000000E0E5D592C000;
defparam prom_inst_0.INIT_RAM_11 = 256'h00008444C00048000000000000000C000000C00000000C000000084444448000;
defparam prom_inst_0.INIT_RAM_12 = 256'h000044480008440000008444444444000000000000000000000044444C444400;
defparam prom_inst_0.INIT_RAM_13 = 256'h0000844444444800000044444C44440000002222222A62000000C00000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h000084448000480000004444884448000004CC44444448000000000008444800;
defparam prom_inst_0.INIT_RAM_15 = 256'h000026A222222200000000884422220000008444444444000000000000000E00;
defparam prom_inst_0.INIT_RAM_16 = 256'h00000000000000000000C00000844C0000000000084422000000444800844400;
defparam prom_inst_0.INIT_RAM_17 = 256'h00C0000000000000000000000000800000000000000000000000880000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h000084000480000000008444448000000000C444C48000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h08444C444480000000000000000048000000840C448000000000C44444C44400;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000448084400000008888888880800000000000000000000000444444800000;
defparam prom_inst_0.INIT_RAM_1B = 256'h000084444480000000004444448000000000222222C000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h000084480480000000000000008000000444C44444C000000000844444800000;
defparam prom_inst_0.INIT_RAM_1D = 256'h00004A222220000000000884422000000000C444444000000000800000800000;
defparam prom_inst_0.INIT_RAM_1E = 256'h00080000000008000000C00008C0000000844C44444000000000248084200000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0006444000000000000000000000840000000000800000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_08 = 256'h000044F444F4400000000000000AAA0000008808888888000000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h0000000000084400000078885344430000000842104AA4000002788007888720;
defparam prom_inst_1.INIT_RAM_0A = 256'h00000022F220000000000043F340000000084222222248000002488888884200;
defparam prom_inst_1.INIT_RAM_0B = 256'h0000884422110000000088000000000000000000F00000000008440000000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h00007800030087000000F884210087000000111111953100000078CAA9988700;
defparam prom_inst_1.INIT_RAM_0D = 256'h0000222210000F00000078888F884300000078000F888F0000000000F8421000;
defparam prom_inst_1.INIT_RAM_0E = 256'h0008440004400000000088000880000000007800078887000000788887888700;
defparam prom_inst_1.INIT_RAM_0F = 256'h000022021008870000008421012480000000000F0F0000000000012484210000;
defparam prom_inst_1.INIT_RAM_10 = 256'h00007888888887000000F8888F888F0000008888F88887000000349A98943000;
defparam prom_inst_1.INIT_RAM_11 = 256'h0000788898888700000088888F888F000000F8888F888F000000F88888888F00;
defparam prom_inst_1.INIT_RAM_12 = 256'h000088889E98880000007880000000000000888888888800000088888F888800;
defparam prom_inst_1.INIT_RAM_13 = 256'h000078888888870000008888889AC80000008888899AC8000000F88888888800;
defparam prom_inst_1.INIT_RAM_14 = 256'h0000780003488700000088888F888F000000789888888700000088888F888F00;
defparam prom_inst_1.INIT_RAM_15 = 256'h00008CA999888800000011224488880000007888888888000000111111111F00;
defparam prom_inst_1.INIT_RAM_16 = 256'h000E888888888E000000F88421000F0000001111124488000000888433488800;
defparam prom_inst_1.INIT_RAM_17 = 256'h00F00000000000000000000000008520000E222222222E000000001122448800;
defparam prom_inst_1.INIT_RAM_18 = 256'h00007888887000000000F88888F8880000007888707000000000000000048800;
defparam prom_inst_1.INIT_RAM_19 = 256'h0780788888700000000044444F4443000000788F887000000000788888700000;
defparam prom_inst_1.INIT_RAM_1A = 256'h0000888F88888800078800000000000000008888888080000000888888F88800;
defparam prom_inst_1.INIT_RAM_1B = 256'h00007888887000000000888888F000000000899999E000000000488888888800;
defparam prom_inst_1.INIT_RAM_1C = 256'h0000780788700000000088888CB0000000007888887000000888F88888F00000;
defparam prom_inst_1.INIT_RAM_1D = 256'h00004A9998800000000012244880000000007888888000000000122222F22000;
defparam prom_inst_1.INIT_RAM_1E = 256'h00012222C22221000000F84210F000000F007888888000000000842124800000;
defparam prom_inst_1.INIT_RAM_1F = 256'h00000032330CAAC00000000000009600000C222212222C000000888880888800;

endmodule //Gowin_pROM_font
