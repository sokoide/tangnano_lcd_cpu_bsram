542: begin adb <= 8'h30; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
544: begin v_ada <= 544; v_din <= to_hexchar(dout[7:4]); end
545: begin v_ada <= 545; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h31; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
546: begin v_ada <= 546; v_din <= to_hexchar(dout[7:4]); end
547: begin v_ada <= 547; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h32; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
548: begin v_ada <= 548; v_din <= to_hexchar(dout[7:4]); end
549: begin v_ada <= 549; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h33; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
550: begin v_ada <= 550; v_din <= to_hexchar(dout[7:4]); end
551: begin v_ada <= 551; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h34; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
553: begin v_ada <= 553; v_din <= to_hexchar(dout[7:4]); end
554: begin v_ada <= 554; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h35; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
555: begin v_ada <= 555; v_din <= to_hexchar(dout[7:4]); end
556: begin v_ada <= 556; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h36; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
557: begin v_ada <= 557; v_din <= to_hexchar(dout[7:4]); end
558: begin v_ada <= 558; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h37; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
559: begin v_ada <= 559; v_din <= to_hexchar(dout[7:4]); end
560: begin v_ada <= 560; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h38; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
563: begin v_ada <= 563; v_din <= to_hexchar(dout[7:4]); end
564: begin v_ada <= 564; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h39; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
565: begin v_ada <= 565; v_din <= to_hexchar(dout[7:4]); end
566: begin v_ada <= 566; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h3A; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
567: begin v_ada <= 567; v_din <= to_hexchar(dout[7:4]); end
568: begin v_ada <= 568; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h3B; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
569: begin v_ada <= 569; v_din <= to_hexchar(dout[7:4]); end
570: begin v_ada <= 570; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h3C; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
572: begin v_ada <= 572; v_din <= to_hexchar(dout[7:4]); end
573: begin v_ada <= 573; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h3D; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
574: begin v_ada <= 574; v_din <= to_hexchar(dout[7:4]); end
575: begin v_ada <= 575; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h3E; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
576: begin v_ada <= 576; v_din <= to_hexchar(dout[7:4]); end
577: begin v_ada <= 577; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h3F; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
578: begin v_ada <= 578; v_din <= to_hexchar(dout[7:4]); end
579: begin v_ada <= 579; v_din <= to_hexchar(dout[3:0]); end
