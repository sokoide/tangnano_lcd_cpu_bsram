422: begin adb <= 8'h10; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
424: begin v_ada <= 424; v_din <= to_hexchar(dout[7:4]); end
425: begin v_ada <= 425; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h11; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
426: begin v_ada <= 426; v_din <= to_hexchar(dout[7:4]); end
427: begin v_ada <= 427; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h12; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
428: begin v_ada <= 428; v_din <= to_hexchar(dout[7:4]); end
429: begin v_ada <= 429; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h13; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
430: begin v_ada <= 430; v_din <= to_hexchar(dout[7:4]); end
431: begin v_ada <= 431; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h14; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
433: begin v_ada <= 433; v_din <= to_hexchar(dout[7:4]); end
434: begin v_ada <= 434; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h15; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
435: begin v_ada <= 435; v_din <= to_hexchar(dout[7:4]); end
436: begin v_ada <= 436; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h16; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
437: begin v_ada <= 437; v_din <= to_hexchar(dout[7:4]); end
438: begin v_ada <= 438; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h17; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
439: begin v_ada <= 439; v_din <= to_hexchar(dout[7:4]); end
440: begin v_ada <= 440; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h18; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
443: begin v_ada <= 443; v_din <= to_hexchar(dout[7:4]); end
444: begin v_ada <= 444; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h19; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
445: begin v_ada <= 445; v_din <= to_hexchar(dout[7:4]); end
446: begin v_ada <= 446; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h1A; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
447: begin v_ada <= 447; v_din <= to_hexchar(dout[7:4]); end
448: begin v_ada <= 448; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h1B; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
449: begin v_ada <= 449; v_din <= to_hexchar(dout[7:4]); end
450: begin v_ada <= 450; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h1C; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
452: begin v_ada <= 452; v_din <= to_hexchar(dout[7:4]); end
453: begin v_ada <= 453; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h1D; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
454: begin v_ada <= 454; v_din <= to_hexchar(dout[7:4]); end
455: begin v_ada <= 455; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h1E; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
456: begin v_ada <= 456; v_din <= to_hexchar(dout[7:4]); end
457: begin v_ada <= 457; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h1F; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
458: begin v_ada <= 458; v_din <= to_hexchar(dout[7:4]); end
459: begin v_ada <= 459; v_din <= to_hexchar(dout[3:0]); end
