602: begin adb <= 8'h40; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
604: begin v_ada <= 604; v_din <= to_hexchar(dout[7:4]); end
605: begin v_ada <= 605; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h41; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
606: begin v_ada <= 606; v_din <= to_hexchar(dout[7:4]); end
607: begin v_ada <= 607; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h42; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
608: begin v_ada <= 608; v_din <= to_hexchar(dout[7:4]); end
609: begin v_ada <= 609; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h43; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
610: begin v_ada <= 610; v_din <= to_hexchar(dout[7:4]); end
611: begin v_ada <= 611; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h44; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
613: begin v_ada <= 613; v_din <= to_hexchar(dout[7:4]); end
614: begin v_ada <= 614; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h45; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
615: begin v_ada <= 615; v_din <= to_hexchar(dout[7:4]); end
616: begin v_ada <= 616; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h46; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
617: begin v_ada <= 617; v_din <= to_hexchar(dout[7:4]); end
618: begin v_ada <= 618; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h47; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
619: begin v_ada <= 619; v_din <= to_hexchar(dout[7:4]); end
620: begin v_ada <= 620; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h48; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
623: begin v_ada <= 623; v_din <= to_hexchar(dout[7:4]); end
624: begin v_ada <= 624; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h49; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
625: begin v_ada <= 625; v_din <= to_hexchar(dout[7:4]); end
626: begin v_ada <= 626; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h4A; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
627: begin v_ada <= 627; v_din <= to_hexchar(dout[7:4]); end
628: begin v_ada <= 628; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h4B; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
629: begin v_ada <= 629; v_din <= to_hexchar(dout[7:4]); end
630: begin v_ada <= 630; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h4C; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
632: begin v_ada <= 632; v_din <= to_hexchar(dout[7:4]); end
633: begin v_ada <= 633; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h4D; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
634: begin v_ada <= 634; v_din <= to_hexchar(dout[7:4]); end
635: begin v_ada <= 635; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h4E; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
636: begin v_ada <= 636; v_din <= to_hexchar(dout[7:4]); end
637: begin v_ada <= 637; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h4F; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z04; end
638: begin v_ada <= 638; v_din <= to_hexchar(dout[7:4]); end
639: begin v_ada <= 639; v_din <= to_hexchar(dout[3:0]); end
