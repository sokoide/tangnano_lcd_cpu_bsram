362: begin adb <= 8'h00; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
364: begin v_ada <= 364; v_din <= to_hexchar(dout[7:4]); end
365: begin v_ada <= 365; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h01; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
366: begin v_ada <= 366; v_din <= to_hexchar(dout[7:4]); end
367: begin v_ada <= 367; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h02; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
368: begin v_ada <= 368; v_din <= to_hexchar(dout[7:4]); end
369: begin v_ada <= 369; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h03; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
370: begin v_ada <= 370; v_din <= to_hexchar(dout[7:4]); end
371: begin v_ada <= 371; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h04; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
373: begin v_ada <= 373; v_din <= to_hexchar(dout[7:4]); end
374: begin v_ada <= 374; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h05; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
375: begin v_ada <= 375; v_din <= to_hexchar(dout[7:4]); end
376: begin v_ada <= 376; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h06; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
377: begin v_ada <= 377; v_din <= to_hexchar(dout[7:4]); end
378: begin v_ada <= 378; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h07; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
379: begin v_ada <= 379; v_din <= to_hexchar(dout[7:4]); end
380: begin v_ada <= 380; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h08; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
383: begin v_ada <= 383; v_din <= to_hexchar(dout[7:4]); end
384: begin v_ada <= 384; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h09; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
385: begin v_ada <= 385; v_din <= to_hexchar(dout[7:4]); end
386: begin v_ada <= 386; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h0A; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
387: begin v_ada <= 387; v_din <= to_hexchar(dout[7:4]); end
388: begin v_ada <= 388; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h0B; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
389: begin v_ada <= 389; v_din <= to_hexchar(dout[7:4]); end
390: begin v_ada <= 390; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h0C; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
392: begin v_ada <= 392; v_din <= to_hexchar(dout[7:4]); end
393: begin v_ada <= 393; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h0D; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
394: begin v_ada <= 394; v_din <= to_hexchar(dout[7:4]); end
395: begin v_ada <= 395; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h0E; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
396: begin v_ada <= 396; v_din <= to_hexchar(dout[7:4]); end
397: begin v_ada <= 397; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h0F; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
398: begin v_ada <= 398; v_din <= to_hexchar(dout[7:4]); end
399: begin v_ada <= 399; v_din <= to_hexchar(dout[3:0]); end
