logic [7:0] boot_program[256];

assign boot_program = '{
        0: 8'hA9,
        1: 8'h41,
        2: 8'h85,
        3: 8'h01,
        4: 8'h8D,
        5: 8'h00,
        6: 8'hE0,
        7: 8'hFF,
        8: 8'h1D,
        9: 8'hDF,
        10: 8'h00,
        11: 8'h00,
        12: 8'hFF,
        13: 8'h1D,
        14: 8'hCF,
        15: 8'h18,
        16: 8'h69,
        17: 8'h01,
        18: 8'hC9,
        19: 8'h46,
        20: 8'hD0,
        21: 8'hEC,
        22: 8'hA9,
        23: 8'h41,
        24: 8'h4C,
        25: 8'h02,
        26: 8'h02,
        default: 8'hEA
    };
parameter logic[7:0] boot_program_length = 27;
