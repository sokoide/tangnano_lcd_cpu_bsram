782: begin adb <= 8'h70; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
784: begin v_ada <= 784; v_din <= to_hexchar(dout[7:4]); end
785: begin v_ada <= 785; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h71; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
786: begin v_ada <= 786; v_din <= to_hexchar(dout[7:4]); end
787: begin v_ada <= 787; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h72; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
788: begin v_ada <= 788; v_din <= to_hexchar(dout[7:4]); end
789: begin v_ada <= 789; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h73; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
790: begin v_ada <= 790; v_din <= to_hexchar(dout[7:4]); end
791: begin v_ada <= 791; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h74; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
793: begin v_ada <= 793; v_din <= to_hexchar(dout[7:4]); end
794: begin v_ada <= 794; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h75; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
795: begin v_ada <= 795; v_din <= to_hexchar(dout[7:4]); end
796: begin v_ada <= 796; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h76; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
797: begin v_ada <= 797; v_din <= to_hexchar(dout[7:4]); end
798: begin v_ada <= 798; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h77; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
799: begin v_ada <= 799; v_din <= to_hexchar(dout[7:4]); end
800: begin v_ada <= 800; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h78; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
803: begin v_ada <= 803; v_din <= to_hexchar(dout[7:4]); end
804: begin v_ada <= 804; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h79; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
805: begin v_ada <= 805; v_din <= to_hexchar(dout[7:4]); end
806: begin v_ada <= 806; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h7A; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
807: begin v_ada <= 807; v_din <= to_hexchar(dout[7:4]); end
808: begin v_ada <= 808; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h7B; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
809: begin v_ada <= 809; v_din <= to_hexchar(dout[7:4]); end
810: begin v_ada <= 810; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h7C; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
812: begin v_ada <= 812; v_din <= to_hexchar(dout[7:4]); end
813: begin v_ada <= 813; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h7D; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
814: begin v_ada <= 814; v_din <= to_hexchar(dout[7:4]); end
815: begin v_ada <= 815; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h7E; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
816: begin v_ada <= 816; v_din <= to_hexchar(dout[7:4]); end
817: begin v_ada <= 817; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h7F; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
818: begin v_ada <= 818; v_din <= to_hexchar(dout[7:4]); end
819: begin v_ada <= 819; v_din <= to_hexchar(dout[3:0]); end
