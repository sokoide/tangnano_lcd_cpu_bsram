722: begin adb <= operands[15:0] + 8'h30 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
724: begin v_ada <= 724; v_din <= to_hexchar(dout[7:4]); end
725: begin v_ada <= 725; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h31 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
726: begin v_ada <= 726; v_din <= to_hexchar(dout[7:4]); end
727: begin v_ada <= 727; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h32 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
728: begin v_ada <= 728; v_din <= to_hexchar(dout[7:4]); end
729: begin v_ada <= 729; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h33 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
730: begin v_ada <= 730; v_din <= to_hexchar(dout[7:4]); end
731: begin v_ada <= 731; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h34 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
733: begin v_ada <= 733; v_din <= to_hexchar(dout[7:4]); end
734: begin v_ada <= 734; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h35 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
735: begin v_ada <= 735; v_din <= to_hexchar(dout[7:4]); end
736: begin v_ada <= 736; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h36 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
737: begin v_ada <= 737; v_din <= to_hexchar(dout[7:4]); end
738: begin v_ada <= 738; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h37 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
739: begin v_ada <= 739; v_din <= to_hexchar(dout[7:4]); end
740: begin v_ada <= 740; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h38 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
743: begin v_ada <= 743; v_din <= to_hexchar(dout[7:4]); end
744: begin v_ada <= 744; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h39 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
745: begin v_ada <= 745; v_din <= to_hexchar(dout[7:4]); end
746: begin v_ada <= 746; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h3A & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
747: begin v_ada <= 747; v_din <= to_hexchar(dout[7:4]); end
748: begin v_ada <= 748; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h3B & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
749: begin v_ada <= 749; v_din <= to_hexchar(dout[7:4]); end
750: begin v_ada <= 750; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h3C & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
752: begin v_ada <= 752; v_din <= to_hexchar(dout[7:4]); end
753: begin v_ada <= 753; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h3D & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
754: begin v_ada <= 754; v_din <= to_hexchar(dout[7:4]); end
755: begin v_ada <= 755; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h3E & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
756: begin v_ada <= 756; v_din <= to_hexchar(dout[7:4]); end
757: begin v_ada <= 757; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h3F & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z03; end
758: begin v_ada <= 758; v_din <= to_hexchar(dout[7:4]); end
759: begin v_ada <= 759; v_din <= to_hexchar(dout[3:0]); end
