`include "consts.svh"
module lcd (
    input logic       PixelClk,
    input logic       nRST,
    input logic [7:0] v_dout,
    input logic [7:0] f_dout,

    output logic        LCD_DE,
    output logic [ 4:0] LCD_B,
    output logic [ 5:0] LCD_G,
    output logic [ 4:0] LCD_R,
    output logic [ 9:0] v_adb,
    output logic [11:0] f_ad
);

  // Horizontal and Vertical pixel counters
  logic [15:0] H_PixelCount;
  logic [15:0] V_PixelCount;

  // Sequential logic for pixel counters
  always_ff @(posedge PixelClk or negedge nRST) begin
    if (!nRST) begin
      V_PixelCount <= 16'd0;
      H_PixelCount <= 16'd0;
    end else if (H_PixelCount == PixelForHS) begin
      H_PixelCount <= 16'd0;
      V_PixelCount <= V_PixelCount + 1'b1;
    end else if (V_PixelCount == PixelForVS) begin
      V_PixelCount <= 16'd0;
      H_PixelCount <= 16'd0;
    end else begin
      H_PixelCount <= H_PixelCount + 1'b1;
    end
  end

  // SYNC-DE MODE
  assign LCD_DE = ((H_PixelCount >= H_BackPorch) &&
                   (H_PixelCount < H_PixelValid + H_BackPorch) &&
                   (V_PixelCount >= V_BackPorch) &&
                   (V_PixelCount < V_PixelValid + V_BackPorch)) ? 1'b1 : 1'b0;


  // character display parameters
  localparam NUMBER_WIDTH = 8;
  localparam NUMBER_HEIGHT = 16;

  // simple 8x16 font
  logic [NUMBER_WIDTH-1:0] font[127:0][NUMBER_HEIGHT-1:0];
  always_comb begin
    // char:
    font[0][0] = 8'h0;
    font[0][1] = 8'h0;
    font[0][2] = 8'h0;
    font[0][3] = 8'h0;
    font[0][4] = 8'h0;
    font[0][5] = 8'h0;
    font[0][6] = 8'h0;
    font[0][7] = 8'h0;
    font[0][8] = 8'h0;
    font[0][9] = 8'h0;
    font[0][10] = 8'h0;
    font[0][11] = 8'h0;
    font[0][12] = 8'h0;
    font[0][13] = 8'h0;
    font[0][14] = 8'h0;
    font[0][15] = 8'h0;
    // char: 
    font[1][0] = 8'h0;
    font[1][1] = 8'h0;
    font[1][2] = 8'h0;
    font[1][3] = 8'h0;
    font[1][4] = 8'h0;
    font[1][5] = 8'h0;
    font[1][6] = 8'h0;
    font[1][7] = 8'h0;
    font[1][8] = 8'h0;
    font[1][9] = 8'h0;
    font[1][10] = 8'h0;
    font[1][11] = 8'h0;
    font[1][12] = 8'h0;
    font[1][13] = 8'h0;
    font[1][14] = 8'h0;
    font[1][15] = 8'h0;
    // char: 
    font[2][0] = 8'h0;
    font[2][1] = 8'h0;
    font[2][2] = 8'h0;
    font[2][3] = 8'h0;
    font[2][4] = 8'h0;
    font[2][5] = 8'h0;
    font[2][6] = 8'h0;
    font[2][7] = 8'h0;
    font[2][8] = 8'h0;
    font[2][9] = 8'h0;
    font[2][10] = 8'h0;
    font[2][11] = 8'h0;
    font[2][12] = 8'h0;
    font[2][13] = 8'h0;
    font[2][14] = 8'h0;
    font[2][15] = 8'h0;
    // char: 
    font[3][0] = 8'h0;
    font[3][1] = 8'h0;
    font[3][2] = 8'h0;
    font[3][3] = 8'h0;
    font[3][4] = 8'h0;
    font[3][5] = 8'h0;
    font[3][6] = 8'h0;
    font[3][7] = 8'h0;
    font[3][8] = 8'h0;
    font[3][9] = 8'h0;
    font[3][10] = 8'h0;
    font[3][11] = 8'h0;
    font[3][12] = 8'h0;
    font[3][13] = 8'h0;
    font[3][14] = 8'h0;
    font[3][15] = 8'h0;
    // char: 
    font[4][0] = 8'h0;
    font[4][1] = 8'h0;
    font[4][2] = 8'h0;
    font[4][3] = 8'h0;
    font[4][4] = 8'h0;
    font[4][5] = 8'h0;
    font[4][6] = 8'h0;
    font[4][7] = 8'h0;
    font[4][8] = 8'h0;
    font[4][9] = 8'h0;
    font[4][10] = 8'h0;
    font[4][11] = 8'h0;
    font[4][12] = 8'h0;
    font[4][13] = 8'h0;
    font[4][14] = 8'h0;
    font[4][15] = 8'h0;
    // char: 
    font[5][0] = 8'h0;
    font[5][1] = 8'h0;
    font[5][2] = 8'h0;
    font[5][3] = 8'h0;
    font[5][4] = 8'h0;
    font[5][5] = 8'h0;
    font[5][6] = 8'h0;
    font[5][7] = 8'h0;
    font[5][8] = 8'h0;
    font[5][9] = 8'h0;
    font[5][10] = 8'h0;
    font[5][11] = 8'h0;
    font[5][12] = 8'h0;
    font[5][13] = 8'h0;
    font[5][14] = 8'h0;
    font[5][15] = 8'h0;
    // char: 
    font[6][0] = 8'h0;
    font[6][1] = 8'h0;
    font[6][2] = 8'h0;
    font[6][3] = 8'h0;
    font[6][4] = 8'h0;
    font[6][5] = 8'h0;
    font[6][6] = 8'h0;
    font[6][7] = 8'h0;
    font[6][8] = 8'h0;
    font[6][9] = 8'h0;
    font[6][10] = 8'h0;
    font[6][11] = 8'h0;
    font[6][12] = 8'h0;
    font[6][13] = 8'h0;
    font[6][14] = 8'h0;
    font[6][15] = 8'h0;
    // char: 
    font[7][0] = 8'h0;
    font[7][1] = 8'h0;
    font[7][2] = 8'h0;
    font[7][3] = 8'h0;
    font[7][4] = 8'h0;
    font[7][5] = 8'h0;
    font[7][6] = 8'h0;
    font[7][7] = 8'h0;
    font[7][8] = 8'h0;
    font[7][9] = 8'h0;
    font[7][10] = 8'h0;
    font[7][11] = 8'h0;
    font[7][12] = 8'h0;
    font[7][13] = 8'h0;
    font[7][14] = 8'h0;
    font[7][15] = 8'h0;
    // char: 
    font[8][0] = 8'h0;
    font[8][1] = 8'h0;
    font[8][2] = 8'h0;
    font[8][3] = 8'h0;
    font[8][4] = 8'h0;
    font[8][5] = 8'h0;
    font[8][6] = 8'h0;
    font[8][7] = 8'h0;
    font[8][8] = 8'h0;
    font[8][9] = 8'h0;
    font[8][10] = 8'h0;
    font[8][11] = 8'h0;
    font[8][12] = 8'h0;
    font[8][13] = 8'h0;
    font[8][14] = 8'h0;
    font[8][15] = 8'h0;
    // char:
    font[9][0] = 8'h0;
    font[9][1] = 8'h0;
    font[9][2] = 8'h0;
    font[9][3] = 8'h0;
    font[9][4] = 8'h0;
    font[9][5] = 8'h0;
    font[9][6] = 8'h0;
    font[9][7] = 8'h0;
    font[9][8] = 8'h0;
    font[9][9] = 8'h0;
    font[9][10] = 8'h0;
    font[9][11] = 8'h0;
    font[9][12] = 8'h0;
    font[9][13] = 8'h0;
    font[9][14] = 8'h0;
    font[9][15] = 8'h0;
    // char:

    font[10][0] = 8'h0;
    font[10][1] = 8'h0;
    font[10][2] = 8'h0;
    font[10][3] = 8'h0;
    font[10][4] = 8'h0;
    font[10][5] = 8'h0;
    font[10][6] = 8'h0;
    font[10][7] = 8'h0;
    font[10][8] = 8'h0;
    font[10][9] = 8'h0;
    font[10][10] = 8'h0;
    font[10][11] = 8'h0;
    font[10][12] = 8'h0;
    font[10][13] = 8'h0;
    font[10][14] = 8'h0;
    font[10][15] = 8'h0;
    // char: 
    font[11][0] = 8'h0;
    font[11][1] = 8'h0;
    font[11][2] = 8'h0;
    font[11][3] = 8'h0;
    font[11][4] = 8'h0;
    font[11][5] = 8'h0;
    font[11][6] = 8'h0;
    font[11][7] = 8'h0;
    font[11][8] = 8'h0;
    font[11][9] = 8'h0;
    font[11][10] = 8'h0;
    font[11][11] = 8'h0;
    font[11][12] = 8'h0;
    font[11][13] = 8'h0;
    font[11][14] = 8'h0;
    font[11][15] = 8'h0;
    // char: 
    font[12][0] = 8'h0;
    font[12][1] = 8'h0;
    font[12][2] = 8'h0;
    font[12][3] = 8'h0;
    font[12][4] = 8'h0;
    font[12][5] = 8'h0;
    font[12][6] = 8'h0;
    font[12][7] = 8'h0;
    font[12][8] = 8'h0;
    font[12][9] = 8'h0;
    font[12][10] = 8'h0;
    font[12][11] = 8'h0;
    font[12][12] = 8'h0;
    font[12][13] = 8'h0;
    font[12][14] = 8'h0;
    font[12][15] = 8'h0;
    // char:
    font[13][0] = 8'h0;
    font[13][1] = 8'h0;
    font[13][2] = 8'h0;
    font[13][3] = 8'h0;
    font[13][4] = 8'h0;
    font[13][5] = 8'h0;
    font[13][6] = 8'h0;
    font[13][7] = 8'h0;
    font[13][8] = 8'h0;
    font[13][9] = 8'h0;
    font[13][10] = 8'h0;
    font[13][11] = 8'h0;
    font[13][12] = 8'h0;
    font[13][13] = 8'h0;
    font[13][14] = 8'h0;
    font[13][15] = 8'h0;
    // char: 
    font[14][0] = 8'h0;
    font[14][1] = 8'h0;
    font[14][2] = 8'h0;
    font[14][3] = 8'h0;
    font[14][4] = 8'h0;
    font[14][5] = 8'h0;
    font[14][6] = 8'h0;
    font[14][7] = 8'h0;
    font[14][8] = 8'h0;
    font[14][9] = 8'h0;
    font[14][10] = 8'h0;
    font[14][11] = 8'h0;
    font[14][12] = 8'h0;
    font[14][13] = 8'h0;
    font[14][14] = 8'h0;
    font[14][15] = 8'h0;
    // char: 
    font[15][0] = 8'h0;
    font[15][1] = 8'h0;
    font[15][2] = 8'h0;
    font[15][3] = 8'h0;
    font[15][4] = 8'h0;
    font[15][5] = 8'h0;
    font[15][6] = 8'h0;
    font[15][7] = 8'h0;
    font[15][8] = 8'h0;
    font[15][9] = 8'h0;
    font[15][10] = 8'h0;
    font[15][11] = 8'h0;
    font[15][12] = 8'h0;
    font[15][13] = 8'h0;
    font[15][14] = 8'h0;
    font[15][15] = 8'h0;
    // char: 
    font[16][0] = 8'h0;
    font[16][1] = 8'h0;
    font[16][2] = 8'h0;
    font[16][3] = 8'h0;
    font[16][4] = 8'h0;
    font[16][5] = 8'h0;
    font[16][6] = 8'h0;
    font[16][7] = 8'h0;
    font[16][8] = 8'h0;
    font[16][9] = 8'h0;
    font[16][10] = 8'h0;
    font[16][11] = 8'h0;
    font[16][12] = 8'h0;
    font[16][13] = 8'h0;
    font[16][14] = 8'h0;
    font[16][15] = 8'h0;
    // char: 
    font[17][0] = 8'h0;
    font[17][1] = 8'h0;
    font[17][2] = 8'h0;
    font[17][3] = 8'h0;
    font[17][4] = 8'h0;
    font[17][5] = 8'h0;
    font[17][6] = 8'h0;
    font[17][7] = 8'h0;
    font[17][8] = 8'h0;
    font[17][9] = 8'h0;
    font[17][10] = 8'h0;
    font[17][11] = 8'h0;
    font[17][12] = 8'h0;
    font[17][13] = 8'h0;
    font[17][14] = 8'h0;
    font[17][15] = 8'h0;
    // char: 
    font[18][0] = 8'h0;
    font[18][1] = 8'h0;
    font[18][2] = 8'h0;
    font[18][3] = 8'h0;
    font[18][4] = 8'h0;
    font[18][5] = 8'h0;
    font[18][6] = 8'h0;
    font[18][7] = 8'h0;
    font[18][8] = 8'h0;
    font[18][9] = 8'h0;
    font[18][10] = 8'h0;
    font[18][11] = 8'h0;
    font[18][12] = 8'h0;
    font[18][13] = 8'h0;
    font[18][14] = 8'h0;
    font[18][15] = 8'h0;
    // char: 
    font[19][0] = 8'h0;
    font[19][1] = 8'h0;
    font[19][2] = 8'h0;
    font[19][3] = 8'h0;
    font[19][4] = 8'h0;
    font[19][5] = 8'h0;
    font[19][6] = 8'h0;
    font[19][7] = 8'h0;
    font[19][8] = 8'h0;
    font[19][9] = 8'h0;
    font[19][10] = 8'h0;
    font[19][11] = 8'h0;
    font[19][12] = 8'h0;
    font[19][13] = 8'h0;
    font[19][14] = 8'h0;
    font[19][15] = 8'h0;
    // char: 
    font[20][0] = 8'h0;
    font[20][1] = 8'h0;
    font[20][2] = 8'h0;
    font[20][3] = 8'h0;
    font[20][4] = 8'h0;
    font[20][5] = 8'h0;
    font[20][6] = 8'h0;
    font[20][7] = 8'h0;
    font[20][8] = 8'h0;
    font[20][9] = 8'h0;
    font[20][10] = 8'h0;
    font[20][11] = 8'h0;
    font[20][12] = 8'h0;
    font[20][13] = 8'h0;
    font[20][14] = 8'h0;
    font[20][15] = 8'h0;
    // char: 
    font[21][0] = 8'h0;
    font[21][1] = 8'h0;
    font[21][2] = 8'h0;
    font[21][3] = 8'h0;
    font[21][4] = 8'h0;
    font[21][5] = 8'h0;
    font[21][6] = 8'h0;
    font[21][7] = 8'h0;
    font[21][8] = 8'h0;
    font[21][9] = 8'h0;
    font[21][10] = 8'h0;
    font[21][11] = 8'h0;
    font[21][12] = 8'h0;
    font[21][13] = 8'h0;
    font[21][14] = 8'h0;
    font[21][15] = 8'h0;
    // char: 
    font[22][0] = 8'h0;
    font[22][1] = 8'h0;
    font[22][2] = 8'h0;
    font[22][3] = 8'h0;
    font[22][4] = 8'h0;
    font[22][5] = 8'h0;
    font[22][6] = 8'h0;
    font[22][7] = 8'h0;
    font[22][8] = 8'h0;
    font[22][9] = 8'h0;
    font[22][10] = 8'h0;
    font[22][11] = 8'h0;
    font[22][12] = 8'h0;
    font[22][13] = 8'h0;
    font[22][14] = 8'h0;
    font[22][15] = 8'h0;
    // char: 
    font[23][0] = 8'h0;
    font[23][1] = 8'h0;
    font[23][2] = 8'h0;
    font[23][3] = 8'h0;
    font[23][4] = 8'h0;
    font[23][5] = 8'h0;
    font[23][6] = 8'h0;
    font[23][7] = 8'h0;
    font[23][8] = 8'h0;
    font[23][9] = 8'h0;
    font[23][10] = 8'h0;
    font[23][11] = 8'h0;
    font[23][12] = 8'h0;
    font[23][13] = 8'h0;
    font[23][14] = 8'h0;
    font[23][15] = 8'h0;
    // char: 
    font[24][0] = 8'h0;
    font[24][1] = 8'h0;
    font[24][2] = 8'h0;
    font[24][3] = 8'h0;
    font[24][4] = 8'h0;
    font[24][5] = 8'h0;
    font[24][6] = 8'h0;
    font[24][7] = 8'h0;
    font[24][8] = 8'h0;
    font[24][9] = 8'h0;
    font[24][10] = 8'h0;
    font[24][11] = 8'h0;
    font[24][12] = 8'h0;
    font[24][13] = 8'h0;
    font[24][14] = 8'h0;
    font[24][15] = 8'h0;
    // char: 
    font[25][0] = 8'h0;
    font[25][1] = 8'h0;
    font[25][2] = 8'h0;
    font[25][3] = 8'h0;
    font[25][4] = 8'h0;
    font[25][5] = 8'h0;
    font[25][6] = 8'h0;
    font[25][7] = 8'h0;
    font[25][8] = 8'h0;
    font[25][9] = 8'h0;
    font[25][10] = 8'h0;
    font[25][11] = 8'h0;
    font[25][12] = 8'h0;
    font[25][13] = 8'h0;
    font[25][14] = 8'h0;
    font[25][15] = 8'h0;
    // char: 
    font[26][0] = 8'h0;
    font[26][1] = 8'h0;
    font[26][2] = 8'h0;
    font[26][3] = 8'h0;
    font[26][4] = 8'h0;
    font[26][5] = 8'h0;
    font[26][6] = 8'h0;
    font[26][7] = 8'h0;
    font[26][8] = 8'h0;
    font[26][9] = 8'h0;
    font[26][10] = 8'h0;
    font[26][11] = 8'h0;
    font[26][12] = 8'h0;
    font[26][13] = 8'h0;
    font[26][14] = 8'h0;
    font[26][15] = 8'h0;
    // char: 
    font[27][0] = 8'h0;
    font[27][1] = 8'h0;
    font[27][2] = 8'h0;
    font[27][3] = 8'h0;
    font[27][4] = 8'h0;
    font[27][5] = 8'h0;
    font[27][6] = 8'h0;
    font[27][7] = 8'h0;
    font[27][8] = 8'h0;
    font[27][9] = 8'h0;
    font[27][10] = 8'h0;
    font[27][11] = 8'h0;
    font[27][12] = 8'h0;
    font[27][13] = 8'h0;
    font[27][14] = 8'h0;
    font[27][15] = 8'h0;
    // char: 
    font[28][0] = 8'h0;
    font[28][1] = 8'h0;
    font[28][2] = 8'h0;
    font[28][3] = 8'h0;
    font[28][4] = 8'h0;
    font[28][5] = 8'h0;
    font[28][6] = 8'h0;
    font[28][7] = 8'h0;
    font[28][8] = 8'h0;
    font[28][9] = 8'h0;
    font[28][10] = 8'h0;
    font[28][11] = 8'h0;
    font[28][12] = 8'h0;
    font[28][13] = 8'h0;
    font[28][14] = 8'h0;
    font[28][15] = 8'h0;
    // char: 
    font[29][0] = 8'h0;
    font[29][1] = 8'h0;
    font[29][2] = 8'h0;
    font[29][3] = 8'h0;
    font[29][4] = 8'h0;
    font[29][5] = 8'h0;
    font[29][6] = 8'h0;
    font[29][7] = 8'h0;
    font[29][8] = 8'h0;
    font[29][9] = 8'h0;
    font[29][10] = 8'h0;
    font[29][11] = 8'h0;
    font[29][12] = 8'h0;
    font[29][13] = 8'h0;
    font[29][14] = 8'h0;
    font[29][15] = 8'h0;
    // char: 
    font[30][0] = 8'h0;
    font[30][1] = 8'h0;
    font[30][2] = 8'h0;
    font[30][3] = 8'h0;
    font[30][4] = 8'h0;
    font[30][5] = 8'h0;
    font[30][6] = 8'h0;
    font[30][7] = 8'h0;
    font[30][8] = 8'h0;
    font[30][9] = 8'h0;
    font[30][10] = 8'h0;
    font[30][11] = 8'h0;
    font[30][12] = 8'h0;
    font[30][13] = 8'h0;
    font[30][14] = 8'h0;
    font[30][15] = 8'h0;
    // char: 
    font[31][0] = 8'h0;
    font[31][1] = 8'h0;
    font[31][2] = 8'h0;
    font[31][3] = 8'h0;
    font[31][4] = 8'h0;
    font[31][5] = 8'h0;
    font[31][6] = 8'h0;
    font[31][7] = 8'h0;
    font[31][8] = 8'h0;
    font[31][9] = 8'h0;
    font[31][10] = 8'h0;
    font[31][11] = 8'h0;
    font[31][12] = 8'h0;
    font[31][13] = 8'h0;
    font[31][14] = 8'h0;
    font[31][15] = 8'h0;
    // char:
    font[32][0] = 8'h0;
    font[32][1] = 8'h0;
    font[32][2] = 8'h0;
    font[32][3] = 8'h0;
    font[32][4] = 8'h0;
    font[32][5] = 8'h0;
    font[32][6] = 8'h0;
    font[32][7] = 8'h0;
    font[32][8] = 8'h0;
    font[32][9] = 8'h0;
    font[32][10] = 8'h0;
    font[32][11] = 8'h0;
    font[32][12] = 8'h0;
    font[32][13] = 8'h0;
    font[32][14] = 8'h0;
    font[32][15] = 8'h0;
    // char: !
    font[33][0] = 8'h0;
    font[33][1] = 8'h0;
    font[33][2] = 8'h80;
    font[33][3] = 8'h80;
    font[33][4] = 8'h80;
    font[33][5] = 8'h80;
    font[33][6] = 8'h80;
    font[33][7] = 8'h80;
    font[33][8] = 8'h80;
    font[33][9] = 8'h0;
    font[33][10] = 8'h80;
    font[33][11] = 8'h80;
    font[33][12] = 8'h0;
    font[33][13] = 8'h0;
    font[33][14] = 8'h0;
    font[33][15] = 8'h0;
    // char: "
    font[34][0] = 8'h0;
    font[34][1] = 8'h0;
    font[34][2] = 8'ha0;
    font[34][3] = 8'ha0;
    font[34][4] = 8'ha0;
    font[34][5] = 8'h0;
    font[34][6] = 8'h0;
    font[34][7] = 8'h0;
    font[34][8] = 8'h0;
    font[34][9] = 8'h0;
    font[34][10] = 8'h0;
    font[34][11] = 8'h0;
    font[34][12] = 8'h0;
    font[34][13] = 8'h0;
    font[34][14] = 8'h0;
    font[34][15] = 8'h0;
    // char: #
    font[35][0] = 8'h0;
    font[35][1] = 8'h0;
    font[35][2] = 8'h0;
    font[35][3] = 8'h48;
    font[35][4] = 8'h48;
    font[35][5] = 8'hfc;
    font[35][6] = 8'h48;
    font[35][7] = 8'h48;
    font[35][8] = 8'h48;
    font[35][9] = 8'hfc;
    font[35][10] = 8'h48;
    font[35][11] = 8'h48;
    font[35][12] = 8'h0;
    font[35][13] = 8'h0;
    font[35][14] = 8'h0;
    font[35][15] = 8'h0;
    // char: $
    font[36][0] = 8'h0;
    font[36][1] = 8'h20;
    font[36][2] = 8'h70;
    font[36][3] = 8'h88;
    font[36][4] = 8'h88;
    font[36][5] = 8'h80;
    font[36][6] = 8'h70;
    font[36][7] = 8'h8;
    font[36][8] = 8'h8;
    font[36][9] = 8'h88;
    font[36][10] = 8'h88;
    font[36][11] = 8'h70;
    font[36][12] = 8'h20;
    font[36][13] = 8'h0;
    font[36][14] = 8'h0;
    font[36][15] = 8'h0;
    // char: %
    font[37][0] = 8'h0;
    font[37][1] = 8'h0;
    font[37][2] = 8'h40;
    font[37][3] = 8'ha0;
    font[37][4] = 8'ha2;
    font[37][5] = 8'h44;
    font[37][6] = 8'h8;
    font[37][7] = 8'h10;
    font[37][8] = 8'h20;
    font[37][9] = 8'h44;
    font[37][10] = 8'h8a;
    font[37][11] = 8'ha;
    font[37][12] = 8'h4;
    font[37][13] = 8'h0;
    font[37][14] = 8'h0;
    font[37][15] = 8'h0;
    // char: &
    font[38][0] = 8'h0;
    font[38][1] = 8'h0;
    font[38][2] = 8'h30;
    font[38][3] = 8'h48;
    font[38][4] = 8'h48;
    font[38][5] = 8'h48;
    font[38][6] = 8'h32;
    font[38][7] = 8'h52;
    font[38][8] = 8'h8c;
    font[38][9] = 8'h84;
    font[38][10] = 8'h8c;
    font[38][11] = 8'h72;
    font[38][12] = 8'h0;
    font[38][13] = 8'h0;
    font[38][14] = 8'h0;
    font[38][15] = 8'h0;
    // char: '
    font[39][0] = 8'h0;
    font[39][1] = 8'h0;
    font[39][2] = 8'h40;
    font[39][3] = 8'h40;
    font[39][4] = 8'h80;
    font[39][5] = 8'h0;
    font[39][6] = 8'h0;
    font[39][7] = 8'h0;
    font[39][8] = 8'h0;
    font[39][9] = 8'h0;
    font[39][10] = 8'h0;
    font[39][11] = 8'h0;
    font[39][12] = 8'h0;
    font[39][13] = 8'h0;
    font[39][14] = 8'h0;
    font[39][15] = 8'h0;
    // char: (
    font[40][0] = 8'h0;
    font[40][1] = 8'h0;
    font[40][2] = 8'h20;
    font[40][3] = 8'h40;
    font[40][4] = 8'h80;
    font[40][5] = 8'h80;
    font[40][6] = 8'h80;
    font[40][7] = 8'h80;
    font[40][8] = 8'h80;
    font[40][9] = 8'h80;
    font[40][10] = 8'h80;
    font[40][11] = 8'h40;
    font[40][12] = 8'h20;
    font[40][13] = 8'h0;
    font[40][14] = 8'h0;
    font[40][15] = 8'h0;
    // char: )
    font[41][0] = 8'h0;
    font[41][1] = 8'h0;
    font[41][2] = 8'h80;
    font[41][3] = 8'h40;
    font[41][4] = 8'h20;
    font[41][5] = 8'h20;
    font[41][6] = 8'h20;
    font[41][7] = 8'h20;
    font[41][8] = 8'h20;
    font[41][9] = 8'h20;
    font[41][10] = 8'h20;
    font[41][11] = 8'h40;
    font[41][12] = 8'h80;
    font[41][13] = 8'h0;
    font[41][14] = 8'h0;
    font[41][15] = 8'h0;
    // char: *
    font[42][0] = 8'h0;
    font[42][1] = 8'h0;
    font[42][2] = 8'h0;
    font[42][3] = 8'h0;
    font[42][4] = 8'h0;
    font[42][5] = 8'h48;
    font[42][6] = 8'h30;
    font[42][7] = 8'hfc;
    font[42][8] = 8'h30;
    font[42][9] = 8'h48;
    font[42][10] = 8'h0;
    font[42][11] = 8'h0;
    font[42][12] = 8'h0;
    font[42][13] = 8'h0;
    font[42][14] = 8'h0;
    font[42][15] = 8'h0;
    // char: +
    font[43][0] = 8'h0;
    font[43][1] = 8'h0;
    font[43][2] = 8'h0;
    font[43][3] = 8'h0;
    font[43][4] = 8'h0;
    font[43][5] = 8'h20;
    font[43][6] = 8'h20;
    font[43][7] = 8'hf8;
    font[43][8] = 8'h20;
    font[43][9] = 8'h20;
    font[43][10] = 8'h0;
    font[43][11] = 8'h0;
    font[43][12] = 8'h0;
    font[43][13] = 8'h0;
    font[43][14] = 8'h0;
    font[43][15] = 8'h0;
    // char: ,
    font[44][0] = 8'h0;
    font[44][1] = 8'h0;
    font[44][2] = 8'h0;
    font[44][3] = 8'h0;
    font[44][4] = 8'h0;
    font[44][5] = 8'h0;
    font[44][6] = 8'h0;
    font[44][7] = 8'h0;
    font[44][8] = 8'h0;
    font[44][9] = 8'h0;
    font[44][10] = 8'h40;
    font[44][11] = 8'h40;
    font[44][12] = 8'h80;
    font[44][13] = 8'h0;
    font[44][14] = 8'h0;
    font[44][15] = 8'h0;
    // char: -
    font[45][0] = 8'h0;
    font[45][1] = 8'h0;
    font[45][2] = 8'h0;
    font[45][3] = 8'h0;
    font[45][4] = 8'h0;
    font[45][5] = 8'h0;
    font[45][6] = 8'h0;
    font[45][7] = 8'hf0;
    font[45][8] = 8'h0;
    font[45][9] = 8'h0;
    font[45][10] = 8'h0;
    font[45][11] = 8'h0;
    font[45][12] = 8'h0;
    font[45][13] = 8'h0;
    font[45][14] = 8'h0;
    font[45][15] = 8'h0;
    // char: .
    font[46][0] = 8'h0;
    font[46][1] = 8'h0;
    font[46][2] = 8'h0;
    font[46][3] = 8'h0;
    font[46][4] = 8'h0;
    font[46][5] = 8'h0;
    font[46][6] = 8'h0;
    font[46][7] = 8'h0;
    font[46][8] = 8'h0;
    font[46][9] = 8'h0;
    font[46][10] = 8'h80;
    font[46][11] = 8'h80;
    font[46][12] = 8'h0;
    font[46][13] = 8'h0;
    font[46][14] = 8'h0;
    font[46][15] = 8'h0;
    // char: /
    font[47][0] = 8'h0;
    font[47][1] = 8'h0;
    font[47][2] = 8'h8;
    font[47][3] = 8'h8;
    font[47][4] = 8'h10;
    font[47][5] = 8'h10;
    font[47][6] = 8'h20;
    font[47][7] = 8'h20;
    font[47][8] = 8'h40;
    font[47][9] = 8'h40;
    font[47][10] = 8'h80;
    font[47][11] = 8'h80;
    font[47][12] = 8'h0;
    font[47][13] = 8'h0;
    font[47][14] = 8'h0;
    font[47][15] = 8'h0;
    // char: 0
    font[48][0] = 8'h0;
    font[48][1] = 8'h0;
    font[48][2] = 8'h78;
    font[48][3] = 8'h84;
    font[48][4] = 8'h8c;
    font[48][5] = 8'h94;
    font[48][6] = 8'h94;
    font[48][7] = 8'ha4;
    font[48][8] = 8'ha4;
    font[48][9] = 8'hc4;
    font[48][10] = 8'h84;
    font[48][11] = 8'h78;
    font[48][12] = 8'h0;
    font[48][13] = 8'h0;
    font[48][14] = 8'h0;
    font[48][15] = 8'h0;
    // char: 1
    font[49][0] = 8'h0;
    font[49][1] = 8'h0;
    font[49][2] = 8'h10;
    font[49][3] = 8'h30;
    font[49][4] = 8'h50;
    font[49][5] = 8'h90;
    font[49][6] = 8'h10;
    font[49][7] = 8'h10;
    font[49][8] = 8'h10;
    font[49][9] = 8'h10;
    font[49][10] = 8'h10;
    font[49][11] = 8'h10;
    font[49][12] = 8'h0;
    font[49][13] = 8'h0;
    font[49][14] = 8'h0;
    font[49][15] = 8'h0;
    // char: 2
    font[50][0] = 8'h0;
    font[50][1] = 8'h0;
    font[50][2] = 8'h78;
    font[50][3] = 8'h84;
    font[50][4] = 8'h4;
    font[50][5] = 8'h8;
    font[50][6] = 8'h10;
    font[50][7] = 8'h20;
    font[50][8] = 8'h40;
    font[50][9] = 8'h80;
    font[50][10] = 8'h80;
    font[50][11] = 8'hfc;
    font[50][12] = 8'h0;
    font[50][13] = 8'h0;
    font[50][14] = 8'h0;
    font[50][15] = 8'h0;
    // char: 3
    font[51][0] = 8'h0;
    font[51][1] = 8'h0;
    font[51][2] = 8'h78;
    font[51][3] = 8'h84;
    font[51][4] = 8'h4;
    font[51][5] = 8'h4;
    font[51][6] = 8'h38;
    font[51][7] = 8'h4;
    font[51][8] = 8'h4;
    font[51][9] = 8'h4;
    font[51][10] = 8'h84;
    font[51][11] = 8'h78;
    font[51][12] = 8'h0;
    font[51][13] = 8'h0;
    font[51][14] = 8'h0;
    font[51][15] = 8'h0;
    // char: 4
    font[52][0] = 8'h0;
    font[52][1] = 8'h0;
    font[52][2] = 8'h8;
    font[52][3] = 8'h18;
    font[52][4] = 8'h28;
    font[52][5] = 8'h48;
    font[52][6] = 8'h88;
    font[52][7] = 8'hfc;
    font[52][8] = 8'h8;
    font[52][9] = 8'h8;
    font[52][10] = 8'h8;
    font[52][11] = 8'h8;
    font[52][12] = 8'h0;
    font[52][13] = 8'h0;
    font[52][14] = 8'h0;
    font[52][15] = 8'h0;
    // char: 5
    font[53][0] = 8'h0;
    font[53][1] = 8'h0;
    font[53][2] = 8'hfc;
    font[53][3] = 8'h80;
    font[53][4] = 8'h80;
    font[53][5] = 8'h80;
    font[53][6] = 8'hf8;
    font[53][7] = 8'h4;
    font[53][8] = 8'h4;
    font[53][9] = 8'h4;
    font[53][10] = 8'h84;
    font[53][11] = 8'h78;
    font[53][12] = 8'h0;
    font[53][13] = 8'h0;
    font[53][14] = 8'h0;
    font[53][15] = 8'h0;
    // char: 6
    font[54][0] = 8'h0;
    font[54][1] = 8'h0;
    font[54][2] = 8'h38;
    font[54][3] = 8'h40;
    font[54][4] = 8'h80;
    font[54][5] = 8'h80;
    font[54][6] = 8'hf8;
    font[54][7] = 8'h84;
    font[54][8] = 8'h84;
    font[54][9] = 8'h84;
    font[54][10] = 8'h84;
    font[54][11] = 8'h78;
    font[54][12] = 8'h0;
    font[54][13] = 8'h0;
    font[54][14] = 8'h0;
    font[54][15] = 8'h0;
    // char: 7
    font[55][0] = 8'h0;
    font[55][1] = 8'h0;
    font[55][2] = 8'hfc;
    font[55][3] = 8'h4;
    font[55][4] = 8'h4;
    font[55][5] = 8'h4;
    font[55][6] = 8'h8;
    font[55][7] = 8'h10;
    font[55][8] = 8'h20;
    font[55][9] = 8'h20;
    font[55][10] = 8'h20;
    font[55][11] = 8'h20;
    font[55][12] = 8'h0;
    font[55][13] = 8'h0;
    font[55][14] = 8'h0;
    font[55][15] = 8'h0;
    // char: 8
    font[56][0] = 8'h0;
    font[56][1] = 8'h0;
    font[56][2] = 8'h78;
    font[56][3] = 8'h84;
    font[56][4] = 8'h84;
    font[56][5] = 8'h84;
    font[56][6] = 8'h78;
    font[56][7] = 8'h84;
    font[56][8] = 8'h84;
    font[56][9] = 8'h84;
    font[56][10] = 8'h84;
    font[56][11] = 8'h78;
    font[56][12] = 8'h0;
    font[56][13] = 8'h0;
    font[56][14] = 8'h0;
    font[56][15] = 8'h0;
    // char: 9
    font[57][0] = 8'h0;
    font[57][1] = 8'h0;
    font[57][2] = 8'h78;
    font[57][3] = 8'h84;
    font[57][4] = 8'h84;
    font[57][5] = 8'h84;
    font[57][6] = 8'h7c;
    font[57][7] = 8'h4;
    font[57][8] = 8'h4;
    font[57][9] = 8'h4;
    font[57][10] = 8'h84;
    font[57][11] = 8'h78;
    font[57][12] = 8'h0;
    font[57][13] = 8'h0;
    font[57][14] = 8'h0;
    font[57][15] = 8'h0;
    // char: :
    font[58][0] = 8'h0;
    font[58][1] = 8'h0;
    font[58][2] = 8'h0;
    font[58][3] = 8'h0;
    font[58][4] = 8'h0;
    font[58][5] = 8'h80;
    font[58][6] = 8'h80;
    font[58][7] = 8'h0;
    font[58][8] = 8'h0;
    font[58][9] = 8'h0;
    font[58][10] = 8'h80;
    font[58][11] = 8'h80;
    font[58][12] = 8'h0;
    font[58][13] = 8'h0;
    font[58][14] = 8'h0;
    font[58][15] = 8'h0;
    // char: ;
    font[59][0] = 8'h0;
    font[59][1] = 8'h0;
    font[59][2] = 8'h0;
    font[59][3] = 8'h0;
    font[59][4] = 8'h0;
    font[59][5] = 8'h40;
    font[59][6] = 8'h40;
    font[59][7] = 8'h0;
    font[59][8] = 8'h0;
    font[59][9] = 8'h0;
    font[59][10] = 8'h40;
    font[59][11] = 8'h40;
    font[59][12] = 8'h80;
    font[59][13] = 8'h0;
    font[59][14] = 8'h0;
    font[59][15] = 8'h0;
    // char: <
    font[60][0] = 8'h0;
    font[60][1] = 8'h0;
    font[60][2] = 8'h0;
    font[60][3] = 8'h8;
    font[60][4] = 8'h10;
    font[60][5] = 8'h20;
    font[60][6] = 8'h40;
    font[60][7] = 8'h80;
    font[60][8] = 8'h40;
    font[60][9] = 8'h20;
    font[60][10] = 8'h10;
    font[60][11] = 8'h8;
    font[60][12] = 8'h0;
    font[60][13] = 8'h0;
    font[60][14] = 8'h0;
    font[60][15] = 8'h0;
    // char: =
    font[61][0] = 8'h0;
    font[61][1] = 8'h0;
    font[61][2] = 8'h0;
    font[61][3] = 8'h0;
    font[61][4] = 8'h0;
    font[61][5] = 8'h0;
    font[61][6] = 8'hfc;
    font[61][7] = 8'h0;
    font[61][8] = 8'hfc;
    font[61][9] = 8'h0;
    font[61][10] = 8'h0;
    font[61][11] = 8'h0;
    font[61][12] = 8'h0;
    font[61][13] = 8'h0;
    font[61][14] = 8'h0;
    font[61][15] = 8'h0;
    // char: >
    font[62][0] = 8'h0;
    font[62][1] = 8'h0;
    font[62][2] = 8'h0;
    font[62][3] = 8'h80;
    font[62][4] = 8'h40;
    font[62][5] = 8'h20;
    font[62][6] = 8'h10;
    font[62][7] = 8'h8;
    font[62][8] = 8'h10;
    font[62][9] = 8'h20;
    font[62][10] = 8'h40;
    font[62][11] = 8'h80;
    font[62][12] = 8'h0;
    font[62][13] = 8'h0;
    font[62][14] = 8'h0;
    font[62][15] = 8'h0;
    // char: ?
    font[63][0] = 8'h0;
    font[63][1] = 8'h0;
    font[63][2] = 8'h78;
    font[63][3] = 8'h84;
    font[63][4] = 8'h84;
    font[63][5] = 8'h4;
    font[63][6] = 8'h8;
    font[63][7] = 8'h10;
    font[63][8] = 8'h20;
    font[63][9] = 8'h0;
    font[63][10] = 8'h20;
    font[63][11] = 8'h20;
    font[63][12] = 8'h0;
    font[63][13] = 8'h0;
    font[63][14] = 8'h0;
    font[63][15] = 8'h0;
    // char: @
    font[64][0] = 8'h0;
    font[64][1] = 8'h0;
    font[64][2] = 8'h0;
    font[64][3] = 8'h3c;
    font[64][4] = 8'h42;
    font[64][5] = 8'h99;
    font[64][6] = 8'h85;
    font[64][7] = 8'h9d;
    font[64][8] = 8'ha5;
    font[64][9] = 8'h9e;
    font[64][10] = 8'h40;
    font[64][11] = 8'h3e;
    font[64][12] = 8'h0;
    font[64][13] = 8'h0;
    font[64][14] = 8'h0;
    font[64][15] = 8'h0;
    // char: A
    font[65][0] = 8'h0;
    font[65][1] = 8'h0;
    font[65][2] = 8'h78;
    font[65][3] = 8'h84;
    font[65][4] = 8'h84;
    font[65][5] = 8'h84;
    font[65][6] = 8'h84;
    font[65][7] = 8'hfc;
    font[65][8] = 8'h84;
    font[65][9] = 8'h84;
    font[65][10] = 8'h84;
    font[65][11] = 8'h84;
    font[65][12] = 8'h0;
    font[65][13] = 8'h0;
    font[65][14] = 8'h0;
    font[65][15] = 8'h0;
    // char: B
    font[66][0] = 8'h0;
    font[66][1] = 8'h0;
    font[66][2] = 8'hf8;
    font[66][3] = 8'h84;
    font[66][4] = 8'h84;
    font[66][5] = 8'h84;
    font[66][6] = 8'hf8;
    font[66][7] = 8'h84;
    font[66][8] = 8'h84;
    font[66][9] = 8'h84;
    font[66][10] = 8'h84;
    font[66][11] = 8'hf8;
    font[66][12] = 8'h0;
    font[66][13] = 8'h0;
    font[66][14] = 8'h0;
    font[66][15] = 8'h0;
    // char: C
    font[67][0] = 8'h0;
    font[67][1] = 8'h0;
    font[67][2] = 8'h78;
    font[67][3] = 8'h84;
    font[67][4] = 8'h80;
    font[67][5] = 8'h80;
    font[67][6] = 8'h80;
    font[67][7] = 8'h80;
    font[67][8] = 8'h80;
    font[67][9] = 8'h80;
    font[67][10] = 8'h84;
    font[67][11] = 8'h78;
    font[67][12] = 8'h0;
    font[67][13] = 8'h0;
    font[67][14] = 8'h0;
    font[67][15] = 8'h0;
    // char: D
    font[68][0] = 8'h0;
    font[68][1] = 8'h0;
    font[68][2] = 8'hf0;
    font[68][3] = 8'h88;
    font[68][4] = 8'h84;
    font[68][5] = 8'h84;
    font[68][6] = 8'h84;
    font[68][7] = 8'h84;
    font[68][8] = 8'h84;
    font[68][9] = 8'h84;
    font[68][10] = 8'h88;
    font[68][11] = 8'hf0;
    font[68][12] = 8'h0;
    font[68][13] = 8'h0;
    font[68][14] = 8'h0;
    font[68][15] = 8'h0;
    // char: E
    font[69][0] = 8'h0;
    font[69][1] = 8'h0;
    font[69][2] = 8'hfc;
    font[69][3] = 8'h80;
    font[69][4] = 8'h80;
    font[69][5] = 8'h80;
    font[69][6] = 8'hf0;
    font[69][7] = 8'h80;
    font[69][8] = 8'h80;
    font[69][9] = 8'h80;
    font[69][10] = 8'h80;
    font[69][11] = 8'hfc;
    font[69][12] = 8'h0;
    font[69][13] = 8'h0;
    font[69][14] = 8'h0;
    font[69][15] = 8'h0;
    // char: F
    font[70][0] = 8'h0;
    font[70][1] = 8'h0;
    font[70][2] = 8'hfc;
    font[70][3] = 8'h80;
    font[70][4] = 8'h80;
    font[70][5] = 8'h80;
    font[70][6] = 8'hf0;
    font[70][7] = 8'h80;
    font[70][8] = 8'h80;
    font[70][9] = 8'h80;
    font[70][10] = 8'h80;
    font[70][11] = 8'h80;
    font[70][12] = 8'h0;
    font[70][13] = 8'h0;
    font[70][14] = 8'h0;
    font[70][15] = 8'h0;
    // char: G
    font[71][0] = 8'h0;
    font[71][1] = 8'h0;
    font[71][2] = 8'h78;
    font[71][3] = 8'h84;
    font[71][4] = 8'h80;
    font[71][5] = 8'h80;
    font[71][6] = 8'h80;
    font[71][7] = 8'h9c;
    font[71][8] = 8'h84;
    font[71][9] = 8'h84;
    font[71][10] = 8'h84;
    font[71][11] = 8'h78;
    font[71][12] = 8'h0;
    font[71][13] = 8'h0;
    font[71][14] = 8'h0;
    font[71][15] = 8'h0;
    // char: H
    font[72][0] = 8'h0;
    font[72][1] = 8'h0;
    font[72][2] = 8'h84;
    font[72][3] = 8'h84;
    font[72][4] = 8'h84;
    font[72][5] = 8'h84;
    font[72][6] = 8'hfc;
    font[72][7] = 8'h84;
    font[72][8] = 8'h84;
    font[72][9] = 8'h84;
    font[72][10] = 8'h84;
    font[72][11] = 8'h84;
    font[72][12] = 8'h0;
    font[72][13] = 8'h0;
    font[72][14] = 8'h0;
    font[72][15] = 8'h0;
    // char: I
    font[73][0] = 8'h0;
    font[73][1] = 8'h0;
    font[73][2] = 8'h80;
    font[73][3] = 8'h80;
    font[73][4] = 8'h80;
    font[73][5] = 8'h80;
    font[73][6] = 8'h80;
    font[73][7] = 8'h80;
    font[73][8] = 8'h80;
    font[73][9] = 8'h80;
    font[73][10] = 8'h80;
    font[73][11] = 8'h80;
    font[73][12] = 8'h0;
    font[73][13] = 8'h0;
    font[73][14] = 8'h0;
    font[73][15] = 8'h0;
    // char: J
    font[74][0] = 8'h0;
    font[74][1] = 8'h0;
    font[74][2] = 8'h4;
    font[74][3] = 8'h4;
    font[74][4] = 8'h4;
    font[74][5] = 8'h4;
    font[74][6] = 8'h4;
    font[74][7] = 8'h4;
    font[74][8] = 8'h4;
    font[74][9] = 8'h84;
    font[74][10] = 8'h84;
    font[74][11] = 8'h78;
    font[74][12] = 8'h0;
    font[74][13] = 8'h0;
    font[74][14] = 8'h0;
    font[74][15] = 8'h0;
    // char: K
    font[75][0] = 8'h0;
    font[75][1] = 8'h0;
    font[75][2] = 8'h84;
    font[75][3] = 8'h84;
    font[75][4] = 8'h88;
    font[75][5] = 8'h90;
    font[75][6] = 8'he0;
    font[75][7] = 8'h90;
    font[75][8] = 8'h88;
    font[75][9] = 8'h84;
    font[75][10] = 8'h84;
    font[75][11] = 8'h84;
    font[75][12] = 8'h0;
    font[75][13] = 8'h0;
    font[75][14] = 8'h0;
    font[75][15] = 8'h0;
    // char: L
    font[76][0] = 8'h0;
    font[76][1] = 8'h0;
    font[76][2] = 8'h80;
    font[76][3] = 8'h80;
    font[76][4] = 8'h80;
    font[76][5] = 8'h80;
    font[76][6] = 8'h80;
    font[76][7] = 8'h80;
    font[76][8] = 8'h80;
    font[76][9] = 8'h80;
    font[76][10] = 8'h80;
    font[76][11] = 8'hfc;
    font[76][12] = 8'h0;
    font[76][13] = 8'h0;
    font[76][14] = 8'h0;
    font[76][15] = 8'h0;
    // char: M
    font[77][0] = 8'h0;
    font[77][1] = 8'h0;
    font[77][2] = 8'h82;
    font[77][3] = 8'hc6;
    font[77][4] = 8'haa;
    font[77][5] = 8'h92;
    font[77][6] = 8'h92;
    font[77][7] = 8'h82;
    font[77][8] = 8'h82;
    font[77][9] = 8'h82;
    font[77][10] = 8'h82;
    font[77][11] = 8'h82;
    font[77][12] = 8'h0;
    font[77][13] = 8'h0;
    font[77][14] = 8'h0;
    font[77][15] = 8'h0;
    // char: N
    font[78][0] = 8'h0;
    font[78][1] = 8'h0;
    font[78][2] = 8'h84;
    font[78][3] = 8'hc4;
    font[78][4] = 8'ha4;
    font[78][5] = 8'h94;
    font[78][6] = 8'h8c;
    font[78][7] = 8'h84;
    font[78][8] = 8'h84;
    font[78][9] = 8'h84;
    font[78][10] = 8'h84;
    font[78][11] = 8'h84;
    font[78][12] = 8'h0;
    font[78][13] = 8'h0;
    font[78][14] = 8'h0;
    font[78][15] = 8'h0;
    // char: O
    font[79][0] = 8'h0;
    font[79][1] = 8'h0;
    font[79][2] = 8'h78;
    font[79][3] = 8'h84;
    font[79][4] = 8'h84;
    font[79][5] = 8'h84;
    font[79][6] = 8'h84;
    font[79][7] = 8'h84;
    font[79][8] = 8'h84;
    font[79][9] = 8'h84;
    font[79][10] = 8'h84;
    font[79][11] = 8'h78;
    font[79][12] = 8'h0;
    font[79][13] = 8'h0;
    font[79][14] = 8'h0;
    font[79][15] = 8'h0;
    // char: P
    font[80][0] = 8'h0;
    font[80][1] = 8'h0;
    font[80][2] = 8'hf8;
    font[80][3] = 8'h84;
    font[80][4] = 8'h84;
    font[80][5] = 8'h84;
    font[80][6] = 8'hf8;
    font[80][7] = 8'h80;
    font[80][8] = 8'h80;
    font[80][9] = 8'h80;
    font[80][10] = 8'h80;
    font[80][11] = 8'h80;
    font[80][12] = 8'h0;
    font[80][13] = 8'h0;
    font[80][14] = 8'h0;
    font[80][15] = 8'h0;
    // char: Q
    font[81][0] = 8'h0;
    font[81][1] = 8'h0;
    font[81][2] = 8'h78;
    font[81][3] = 8'h84;
    font[81][4] = 8'h84;
    font[81][5] = 8'h84;
    font[81][6] = 8'h84;
    font[81][7] = 8'h84;
    font[81][8] = 8'h84;
    font[81][9] = 8'h94;
    font[81][10] = 8'h8c;
    font[81][11] = 8'h7c;
    font[81][12] = 8'h4;
    font[81][13] = 8'h0;
    font[81][14] = 8'h0;
    font[81][15] = 8'h0;
    // char: R
    font[82][0] = 8'h0;
    font[82][1] = 8'h0;
    font[82][2] = 8'hf8;
    font[82][3] = 8'h84;
    font[82][4] = 8'h84;
    font[82][5] = 8'h84;
    font[82][6] = 8'hf8;
    font[82][7] = 8'h88;
    font[82][8] = 8'h84;
    font[82][9] = 8'h84;
    font[82][10] = 8'h84;
    font[82][11] = 8'h84;
    font[82][12] = 8'h0;
    font[82][13] = 8'h0;
    font[82][14] = 8'h0;
    font[82][15] = 8'h0;
    // char: S
    font[83][0] = 8'h0;
    font[83][1] = 8'h0;
    font[83][2] = 8'h78;
    font[83][3] = 8'h84;
    font[83][4] = 8'h80;
    font[83][5] = 8'h40;
    font[83][6] = 8'h30;
    font[83][7] = 8'h8;
    font[83][8] = 8'h4;
    font[83][9] = 8'h4;
    font[83][10] = 8'h84;
    font[83][11] = 8'h78;
    font[83][12] = 8'h0;
    font[83][13] = 8'h0;
    font[83][14] = 8'h0;
    font[83][15] = 8'h0;
    // char: T
    font[84][0] = 8'h0;
    font[84][1] = 8'h0;
    font[84][2] = 8'hfe;
    font[84][3] = 8'h10;
    font[84][4] = 8'h10;
    font[84][5] = 8'h10;
    font[84][6] = 8'h10;
    font[84][7] = 8'h10;
    font[84][8] = 8'h10;
    font[84][9] = 8'h10;
    font[84][10] = 8'h10;
    font[84][11] = 8'h10;
    font[84][12] = 8'h0;
    font[84][13] = 8'h0;
    font[84][14] = 8'h0;
    font[84][15] = 8'h0;
    // char: U
    font[85][0] = 8'h0;
    font[85][1] = 8'h0;
    font[85][2] = 8'h84;
    font[85][3] = 8'h84;
    font[85][4] = 8'h84;
    font[85][5] = 8'h84;
    font[85][6] = 8'h84;
    font[85][7] = 8'h84;
    font[85][8] = 8'h84;
    font[85][9] = 8'h84;
    font[85][10] = 8'h84;
    font[85][11] = 8'h78;
    font[85][12] = 8'h0;
    font[85][13] = 8'h0;
    font[85][14] = 8'h0;
    font[85][15] = 8'h0;
    // char: V
    font[86][0] = 8'h0;
    font[86][1] = 8'h0;
    font[86][2] = 8'h82;
    font[86][3] = 8'h82;
    font[86][4] = 8'h82;
    font[86][5] = 8'h82;
    font[86][6] = 8'h44;
    font[86][7] = 8'h44;
    font[86][8] = 8'h28;
    font[86][9] = 8'h28;
    font[86][10] = 8'h10;
    font[86][11] = 8'h10;
    font[86][12] = 8'h0;
    font[86][13] = 8'h0;
    font[86][14] = 8'h0;
    font[86][15] = 8'h0;
    // char: W
    font[87][0] = 8'h0;
    font[87][1] = 8'h0;
    font[87][2] = 8'h82;
    font[87][3] = 8'h82;
    font[87][4] = 8'h82;
    font[87][5] = 8'h82;
    font[87][6] = 8'h92;
    font[87][7] = 8'h92;
    font[87][8] = 8'h92;
    font[87][9] = 8'haa;
    font[87][10] = 8'hc6;
    font[87][11] = 8'h82;
    font[87][12] = 8'h0;
    font[87][13] = 8'h0;
    font[87][14] = 8'h0;
    font[87][15] = 8'h0;
    // char: X
    font[88][0] = 8'h0;
    font[88][1] = 8'h0;
    font[88][2] = 8'h84;
    font[88][3] = 8'h84;
    font[88][4] = 8'h84;
    font[88][5] = 8'h48;
    font[88][6] = 8'h30;
    font[88][7] = 8'h30;
    font[88][8] = 8'h48;
    font[88][9] = 8'h84;
    font[88][10] = 8'h84;
    font[88][11] = 8'h84;
    font[88][12] = 8'h0;
    font[88][13] = 8'h0;
    font[88][14] = 8'h0;
    font[88][15] = 8'h0;
    // char: Y
    font[89][0] = 8'h0;
    font[89][1] = 8'h0;
    font[89][2] = 8'h82;
    font[89][3] = 8'h82;
    font[89][4] = 8'h44;
    font[89][5] = 8'h44;
    font[89][6] = 8'h28;
    font[89][7] = 8'h10;
    font[89][8] = 8'h10;
    font[89][9] = 8'h10;
    font[89][10] = 8'h10;
    font[89][11] = 8'h10;
    font[89][12] = 8'h0;
    font[89][13] = 8'h0;
    font[89][14] = 8'h0;
    font[89][15] = 8'h0;
    // char: Z
    font[90][0] = 8'h0;
    font[90][1] = 8'h0;
    font[90][2] = 8'hfc;
    font[90][3] = 8'h4;
    font[90][4] = 8'h4;
    font[90][5] = 8'h8;
    font[90][6] = 8'h10;
    font[90][7] = 8'h20;
    font[90][8] = 8'h40;
    font[90][9] = 8'h80;
    font[90][10] = 8'h80;
    font[90][11] = 8'hfc;
    font[90][12] = 8'h0;
    font[90][13] = 8'h0;
    font[90][14] = 8'h0;
    font[90][15] = 8'h0;
    // char: [
    font[91][0] = 8'h0;
    font[91][1] = 8'h0;
    font[91][2] = 8'he0;
    font[91][3] = 8'h80;
    font[91][4] = 8'h80;
    font[91][5] = 8'h80;
    font[91][6] = 8'h80;
    font[91][7] = 8'h80;
    font[91][8] = 8'h80;
    font[91][9] = 8'h80;
    font[91][10] = 8'h80;
    font[91][11] = 8'h80;
    font[91][12] = 8'he0;
    font[91][13] = 8'h0;
    font[91][14] = 8'h0;
    font[91][15] = 8'h0;
    // char: \
font[92][0] = 8'h0;
    font[92][1] = 8'h0;
    font[92][2] = 8'h80;
    font[92][3] = 8'h80;
    font[92][4] = 8'h40;
    font[92][5] = 8'h40;
    font[92][6] = 8'h20;
    font[92][7] = 8'h20;
    font[92][8] = 8'h10;
    font[92][9] = 8'h10;
    font[92][10] = 8'h8;
    font[92][11] = 8'h8;
    font[92][12] = 8'h0;
    font[92][13] = 8'h0;
    font[92][14] = 8'h0;
    font[92][15] = 8'h0;
    // char: ]
    font[93][0] = 8'h0;
    font[93][1] = 8'h0;
    font[93][2] = 8'he0;
    font[93][3] = 8'h20;
    font[93][4] = 8'h20;
    font[93][5] = 8'h20;
    font[93][6] = 8'h20;
    font[93][7] = 8'h20;
    font[93][8] = 8'h20;
    font[93][9] = 8'h20;
    font[93][10] = 8'h20;
    font[93][11] = 8'h20;
    font[93][12] = 8'he0;
    font[93][13] = 8'h0;
    font[93][14] = 8'h0;
    font[93][15] = 8'h0;
    // char: ^
    font[94][0] = 8'h0;
    font[94][1] = 8'h20;
    font[94][2] = 8'h50;
    font[94][3] = 8'h88;
    font[94][4] = 8'h0;
    font[94][5] = 8'h0;
    font[94][6] = 8'h0;
    font[94][7] = 8'h0;
    font[94][8] = 8'h0;
    font[94][9] = 8'h0;
    font[94][10] = 8'h0;
    font[94][11] = 8'h0;
    font[94][12] = 8'h0;
    font[94][13] = 8'h0;
    font[94][14] = 8'h0;
    font[94][15] = 8'h0;
    // char: _
    font[95][0] = 8'h0;
    font[95][1] = 8'h0;
    font[95][2] = 8'h0;
    font[95][3] = 8'h0;
    font[95][4] = 8'h0;
    font[95][5] = 8'h0;
    font[95][6] = 8'h0;
    font[95][7] = 8'h0;
    font[95][8] = 8'h0;
    font[95][9] = 8'h0;
    font[95][10] = 8'h0;
    font[95][11] = 8'h0;
    font[95][12] = 8'h0;
    font[95][13] = 8'hfc;
    font[95][14] = 8'h0;
    font[95][15] = 8'h0;
    // char: `
    font[96][0] = 8'h0;
    font[96][1] = 8'h0;
    font[96][2] = 8'h80;
    font[96][3] = 8'h80;
    font[96][4] = 8'h40;
    font[96][5] = 8'h0;
    font[96][6] = 8'h0;
    font[96][7] = 8'h0;
    font[96][8] = 8'h0;
    font[96][9] = 8'h0;
    font[96][10] = 8'h0;
    font[96][11] = 8'h0;
    font[96][12] = 8'h0;
    font[96][13] = 8'h0;
    font[96][14] = 8'h0;
    font[96][15] = 8'h0;
    // char: a
    font[97][0] = 8'h0;
    font[97][1] = 8'h0;
    font[97][2] = 8'h0;
    font[97][3] = 8'h0;
    font[97][4] = 8'h0;
    font[97][5] = 8'h78;
    font[97][6] = 8'h4;
    font[97][7] = 8'h7c;
    font[97][8] = 8'h84;
    font[97][9] = 8'h84;
    font[97][10] = 8'h84;
    font[97][11] = 8'h7c;
    font[97][12] = 8'h0;
    font[97][13] = 8'h0;
    font[97][14] = 8'h0;
    font[97][15] = 8'h0;
    // char: b
    font[98][0] = 8'h0;
    font[98][1] = 8'h0;
    font[98][2] = 8'h80;
    font[98][3] = 8'h80;
    font[98][4] = 8'h80;
    font[98][5] = 8'hf8;
    font[98][6] = 8'h84;
    font[98][7] = 8'h84;
    font[98][8] = 8'h84;
    font[98][9] = 8'h84;
    font[98][10] = 8'h84;
    font[98][11] = 8'hf8;
    font[98][12] = 8'h0;
    font[98][13] = 8'h0;
    font[98][14] = 8'h0;
    font[98][15] = 8'h0;
    // char: c
    font[99][0] = 8'h0;
    font[99][1] = 8'h0;
    font[99][2] = 8'h0;
    font[99][3] = 8'h0;
    font[99][4] = 8'h0;
    font[99][5] = 8'h78;
    font[99][6] = 8'h84;
    font[99][7] = 8'h80;
    font[99][8] = 8'h80;
    font[99][9] = 8'h80;
    font[99][10] = 8'h84;
    font[99][11] = 8'h78;
    font[99][12] = 8'h0;
    font[99][13] = 8'h0;
    font[99][14] = 8'h0;
    font[99][15] = 8'h0;
    // char: d
    font[100][0] = 8'h0;
    font[100][1] = 8'h0;
    font[100][2] = 8'h4;
    font[100][3] = 8'h4;
    font[100][4] = 8'h4;
    font[100][5] = 8'h7c;
    font[100][6] = 8'h84;
    font[100][7] = 8'h84;
    font[100][8] = 8'h84;
    font[100][9] = 8'h84;
    font[100][10] = 8'h84;
    font[100][11] = 8'h7c;
    font[100][12] = 8'h0;
    font[100][13] = 8'h0;
    font[100][14] = 8'h0;
    font[100][15] = 8'h0;
    // char: e
    font[101][0] = 8'h0;
    font[101][1] = 8'h0;
    font[101][2] = 8'h0;
    font[101][3] = 8'h0;
    font[101][4] = 8'h0;
    font[101][5] = 8'h78;
    font[101][6] = 8'h84;
    font[101][7] = 8'h84;
    font[101][8] = 8'hfc;
    font[101][9] = 8'h80;
    font[101][10] = 8'h84;
    font[101][11] = 8'h78;
    font[101][12] = 8'h0;
    font[101][13] = 8'h0;
    font[101][14] = 8'h0;
    font[101][15] = 8'h0;
    // char: f
    font[102][0] = 8'h0;
    font[102][1] = 8'h0;
    font[102][2] = 8'h38;
    font[102][3] = 8'h44;
    font[102][4] = 8'h40;
    font[102][5] = 8'h40;
    font[102][6] = 8'hf0;
    font[102][7] = 8'h40;
    font[102][8] = 8'h40;
    font[102][9] = 8'h40;
    font[102][10] = 8'h40;
    font[102][11] = 8'h40;
    font[102][12] = 8'h0;
    font[102][13] = 8'h0;
    font[102][14] = 8'h0;
    font[102][15] = 8'h0;
    // char: g
    font[103][0] = 8'h0;
    font[103][1] = 8'h0;
    font[103][2] = 8'h0;
    font[103][3] = 8'h0;
    font[103][4] = 8'h0;
    font[103][5] = 8'h78;
    font[103][6] = 8'h84;
    font[103][7] = 8'h84;
    font[103][8] = 8'h84;
    font[103][9] = 8'h84;
    font[103][10] = 8'h8c;
    font[103][11] = 8'h74;
    font[103][12] = 8'h4;
    font[103][13] = 8'h84;
    font[103][14] = 8'h78;
    font[103][15] = 8'h0;
    // char: h
    font[104][0] = 8'h0;
    font[104][1] = 8'h0;
    font[104][2] = 8'h80;
    font[104][3] = 8'h80;
    font[104][4] = 8'h80;
    font[104][5] = 8'hf8;
    font[104][6] = 8'h84;
    font[104][7] = 8'h84;
    font[104][8] = 8'h84;
    font[104][9] = 8'h84;
    font[104][10] = 8'h84;
    font[104][11] = 8'h84;
    font[104][12] = 8'h0;
    font[104][13] = 8'h0;
    font[104][14] = 8'h0;
    font[104][15] = 8'h0;
    // char: i
    font[105][0] = 8'h0;
    font[105][1] = 8'h0;
    font[105][2] = 8'h0;
    font[105][3] = 8'h80;
    font[105][4] = 8'h0;
    font[105][5] = 8'h80;
    font[105][6] = 8'h80;
    font[105][7] = 8'h80;
    font[105][8] = 8'h80;
    font[105][9] = 8'h80;
    font[105][10] = 8'h80;
    font[105][11] = 8'h80;
    font[105][12] = 8'h0;
    font[105][13] = 8'h0;
    font[105][14] = 8'h0;
    font[105][15] = 8'h0;
    // char: j
    font[106][0] = 8'h0;
    font[106][1] = 8'h0;
    font[106][2] = 8'h0;
    font[106][3] = 8'h8;
    font[106][4] = 8'h0;
    font[106][5] = 8'h8;
    font[106][6] = 8'h8;
    font[106][7] = 8'h8;
    font[106][8] = 8'h8;
    font[106][9] = 8'h8;
    font[106][10] = 8'h8;
    font[106][11] = 8'h8;
    font[106][12] = 8'h88;
    font[106][13] = 8'h88;
    font[106][14] = 8'h70;
    font[106][15] = 8'h0;
    // char: k
    font[107][0] = 8'h0;
    font[107][1] = 8'h0;
    font[107][2] = 8'h80;
    font[107][3] = 8'h80;
    font[107][4] = 8'h80;
    font[107][5] = 8'h84;
    font[107][6] = 8'h84;
    font[107][7] = 8'h88;
    font[107][8] = 8'hf0;
    font[107][9] = 8'h88;
    font[107][10] = 8'h84;
    font[107][11] = 8'h84;
    font[107][12] = 8'h0;
    font[107][13] = 8'h0;
    font[107][14] = 8'h0;
    font[107][15] = 8'h0;
    // char: l
    font[108][0] = 8'h0;
    font[108][1] = 8'h0;
    font[108][2] = 8'h80;
    font[108][3] = 8'h80;
    font[108][4] = 8'h80;
    font[108][5] = 8'h80;
    font[108][6] = 8'h80;
    font[108][7] = 8'h80;
    font[108][8] = 8'h80;
    font[108][9] = 8'h80;
    font[108][10] = 8'h80;
    font[108][11] = 8'h40;
    font[108][12] = 8'h0;
    font[108][13] = 8'h0;
    font[108][14] = 8'h0;
    font[108][15] = 8'h0;
    // char: m
    font[109][0] = 8'h0;
    font[109][1] = 8'h0;
    font[109][2] = 8'h0;
    font[109][3] = 8'h0;
    font[109][4] = 8'h0;
    font[109][5] = 8'hec;
    font[109][6] = 8'h92;
    font[109][7] = 8'h92;
    font[109][8] = 8'h92;
    font[109][9] = 8'h92;
    font[109][10] = 8'h92;
    font[109][11] = 8'h82;
    font[109][12] = 8'h0;
    font[109][13] = 8'h0;
    font[109][14] = 8'h0;
    font[109][15] = 8'h0;
    // char: n
    font[110][0] = 8'h0;
    font[110][1] = 8'h0;
    font[110][2] = 8'h0;
    font[110][3] = 8'h0;
    font[110][4] = 8'h0;
    font[110][5] = 8'hf8;
    font[110][6] = 8'h84;
    font[110][7] = 8'h84;
    font[110][8] = 8'h84;
    font[110][9] = 8'h84;
    font[110][10] = 8'h84;
    font[110][11] = 8'h84;
    font[110][12] = 8'h0;
    font[110][13] = 8'h0;
    font[110][14] = 8'h0;
    font[110][15] = 8'h0;
    // char: o
    font[111][0] = 8'h0;
    font[111][1] = 8'h0;
    font[111][2] = 8'h0;
    font[111][3] = 8'h0;
    font[111][4] = 8'h0;
    font[111][5] = 8'h78;
    font[111][6] = 8'h84;
    font[111][7] = 8'h84;
    font[111][8] = 8'h84;
    font[111][9] = 8'h84;
    font[111][10] = 8'h84;
    font[111][11] = 8'h78;
    font[111][12] = 8'h0;
    font[111][13] = 8'h0;
    font[111][14] = 8'h0;
    font[111][15] = 8'h0;
    // char: p
    font[112][0] = 8'h0;
    font[112][1] = 8'h0;
    font[112][2] = 8'h0;
    font[112][3] = 8'h0;
    font[112][4] = 8'h0;
    font[112][5] = 8'hf8;
    font[112][6] = 8'h84;
    font[112][7] = 8'h84;
    font[112][8] = 8'h84;
    font[112][9] = 8'h84;
    font[112][10] = 8'h84;
    font[112][11] = 8'hf8;
    font[112][12] = 8'h80;
    font[112][13] = 8'h80;
    font[112][14] = 8'h80;
    font[112][15] = 8'h0;
    // char: q
    font[113][0] = 8'h0;
    font[113][1] = 8'h0;
    font[113][2] = 8'h0;
    font[113][3] = 8'h0;
    font[113][4] = 8'h0;
    font[113][5] = 8'h7c;
    font[113][6] = 8'h84;
    font[113][7] = 8'h84;
    font[113][8] = 8'h84;
    font[113][9] = 8'h84;
    font[113][10] = 8'h84;
    font[113][11] = 8'h7c;
    font[113][12] = 8'h4;
    font[113][13] = 8'h4;
    font[113][14] = 8'h4;
    font[113][15] = 8'h0;
    // char: r
    font[114][0] = 8'h0;
    font[114][1] = 8'h0;
    font[114][2] = 8'h0;
    font[114][3] = 8'h0;
    font[114][4] = 8'h0;
    font[114][5] = 8'hb8;
    font[114][6] = 8'hc0;
    font[114][7] = 8'h80;
    font[114][8] = 8'h80;
    font[114][9] = 8'h80;
    font[114][10] = 8'h80;
    font[114][11] = 8'h80;
    font[114][12] = 8'h0;
    font[114][13] = 8'h0;
    font[114][14] = 8'h0;
    font[114][15] = 8'h0;
    // char: s
    font[115][0] = 8'h0;
    font[115][1] = 8'h0;
    font[115][2] = 8'h0;
    font[115][3] = 8'h0;
    font[115][4] = 8'h0;
    font[115][5] = 8'h78;
    font[115][6] = 8'h84;
    font[115][7] = 8'h80;
    font[115][8] = 8'h78;
    font[115][9] = 8'h4;
    font[115][10] = 8'h84;
    font[115][11] = 8'h78;
    font[115][12] = 8'h0;
    font[115][13] = 8'h0;
    font[115][14] = 8'h0;
    font[115][15] = 8'h0;
    // char: t
    font[116][0] = 8'h0;
    font[116][1] = 8'h0;
    font[116][2] = 8'h0;
    font[116][3] = 8'h20;
    font[116][4] = 8'h20;
    font[116][5] = 8'hf8;
    font[116][6] = 8'h20;
    font[116][7] = 8'h20;
    font[116][8] = 8'h20;
    font[116][9] = 8'h20;
    font[116][10] = 8'h20;
    font[116][11] = 8'h18;
    font[116][12] = 8'h0;
    font[116][13] = 8'h0;
    font[116][14] = 8'h0;
    font[116][15] = 8'h0;
    // char: u
    font[117][0] = 8'h0;
    font[117][1] = 8'h0;
    font[117][2] = 8'h0;
    font[117][3] = 8'h0;
    font[117][4] = 8'h0;
    font[117][5] = 8'h84;
    font[117][6] = 8'h84;
    font[117][7] = 8'h84;
    font[117][8] = 8'h84;
    font[117][9] = 8'h84;
    font[117][10] = 8'h84;
    font[117][11] = 8'h7c;
    font[117][12] = 8'h0;
    font[117][13] = 8'h0;
    font[117][14] = 8'h0;
    font[117][15] = 8'h0;
    // char: v
    font[118][0] = 8'h0;
    font[118][1] = 8'h0;
    font[118][2] = 8'h0;
    font[118][3] = 8'h0;
    font[118][4] = 8'h0;
    font[118][5] = 8'h82;
    font[118][6] = 8'h82;
    font[118][7] = 8'h44;
    font[118][8] = 8'h44;
    font[118][9] = 8'h28;
    font[118][10] = 8'h28;
    font[118][11] = 8'h10;
    font[118][12] = 8'h0;
    font[118][13] = 8'h0;
    font[118][14] = 8'h0;
    font[118][15] = 8'h0;
    // char: w
    font[119][0] = 8'h0;
    font[119][1] = 8'h0;
    font[119][2] = 8'h0;
    font[119][3] = 8'h0;
    font[119][4] = 8'h0;
    font[119][5] = 8'h82;
    font[119][6] = 8'h82;
    font[119][7] = 8'h92;
    font[119][8] = 8'h92;
    font[119][9] = 8'h92;
    font[119][10] = 8'haa;
    font[119][11] = 8'h44;
    font[119][12] = 8'h0;
    font[119][13] = 8'h0;
    font[119][14] = 8'h0;
    font[119][15] = 8'h0;
    // char: x
    font[120][0] = 8'h0;
    font[120][1] = 8'h0;
    font[120][2] = 8'h0;
    font[120][3] = 8'h0;
    font[120][4] = 8'h0;
    font[120][5] = 8'h82;
    font[120][6] = 8'h44;
    font[120][7] = 8'h28;
    font[120][8] = 8'h10;
    font[120][9] = 8'h28;
    font[120][10] = 8'h44;
    font[120][11] = 8'h82;
    font[120][12] = 8'h0;
    font[120][13] = 8'h0;
    font[120][14] = 8'h0;
    font[120][15] = 8'h0;
    // char: y
    font[121][0] = 8'h0;
    font[121][1] = 8'h0;
    font[121][2] = 8'h0;
    font[121][3] = 8'h0;
    font[121][4] = 8'h0;
    font[121][5] = 8'h84;
    font[121][6] = 8'h84;
    font[121][7] = 8'h84;
    font[121][8] = 8'h84;
    font[121][9] = 8'h84;
    font[121][10] = 8'h8c;
    font[121][11] = 8'h74;
    font[121][12] = 8'h4;
    font[121][13] = 8'h8;
    font[121][14] = 8'hf0;
    font[121][15] = 8'h0;
    // char: z
    font[122][0] = 8'h0;
    font[122][1] = 8'h0;
    font[122][2] = 8'h0;
    font[122][3] = 8'h0;
    font[122][4] = 8'h0;
    font[122][5] = 8'hfc;
    font[122][6] = 8'h8;
    font[122][7] = 8'h10;
    font[122][8] = 8'h20;
    font[122][9] = 8'h40;
    font[122][10] = 8'h80;
    font[122][11] = 8'hfc;
    font[122][12] = 8'h0;
    font[122][13] = 8'h0;
    font[122][14] = 8'h0;
    font[122][15] = 8'h0;
    // char: {
    font[123][0] = 8'h0;
    font[123][1] = 8'h0;
    font[123][2] = 8'h18;
    font[123][3] = 8'h20;
    font[123][4] = 8'h20;
    font[123][5] = 8'h20;
    font[123][6] = 8'h20;
    font[123][7] = 8'hc0;
    font[123][8] = 8'h20;
    font[123][9] = 8'h20;
    font[123][10] = 8'h20;
    font[123][11] = 8'h20;
    font[123][12] = 8'h18;
    font[123][13] = 8'h0;
    font[123][14] = 8'h0;
    font[123][15] = 8'h0;
    // char: |
    font[124][0] = 8'h0;
    font[124][1] = 8'h0;
    font[124][2] = 8'h80;
    font[124][3] = 8'h80;
    font[124][4] = 8'h80;
    font[124][5] = 8'h80;
    font[124][6] = 8'h0;
    font[124][7] = 8'h80;
    font[124][8] = 8'h80;
    font[124][9] = 8'h80;
    font[124][10] = 8'h80;
    font[124][11] = 8'h80;
    font[124][12] = 8'h0;
    font[124][13] = 8'h0;
    font[124][14] = 8'h0;
    font[124][15] = 8'h0;
    // char: }
    font[125][0] = 8'h0;
    font[125][1] = 8'h0;
    font[125][2] = 8'hc0;
    font[125][3] = 8'h20;
    font[125][4] = 8'h20;
    font[125][5] = 8'h20;
    font[125][6] = 8'h20;
    font[125][7] = 8'h18;
    font[125][8] = 8'h20;
    font[125][9] = 8'h20;
    font[125][10] = 8'h20;
    font[125][11] = 8'h20;
    font[125][12] = 8'hc0;
    font[125][13] = 8'h0;
    font[125][14] = 8'h0;
    font[125][15] = 8'h0;
    // char: ~
    font[126][0] = 8'h0;
    font[126][1] = 8'h0;
    font[126][2] = 8'h64;
    font[126][3] = 8'h98;
    font[126][4] = 8'h0;
    font[126][5] = 8'h0;
    font[126][6] = 8'h0;
    font[126][7] = 8'h0;
    font[126][8] = 8'h0;
    font[126][9] = 8'h0;
    font[126][10] = 8'h0;
    font[126][11] = 8'h0;
    font[126][12] = 8'h0;
    font[126][13] = 8'h0;
    font[126][14] = 8'h0;
    font[126][15] = 8'h0;
    // char: 
    font[127][0] = 8'h0;
    font[127][1] = 8'hc0;
    font[127][2] = 8'ha0;
    font[127][3] = 8'ha0;
    font[127][4] = 8'hc0;
    font[127][5] = 8'h0;
    font[127][6] = 8'h30;
    font[127][7] = 8'h30;
    font[127][8] = 8'h20;
    font[127][9] = 8'h34;
    font[127][10] = 8'h4;
    font[127][11] = 8'h4;
    font[127][12] = 8'h6;
    font[127][13] = 8'h0;
    font[127][14] = 8'h0;
    font[127][15] = 8'h0;
  end


  logic [7:0] char;

  always_ff @(posedge PixelClk or negedge nRST) begin
    // x could be minus (underflow) when H_PixelCount is smaller than H_BackPorch
    // so we need to use signed logic to avoid the underflow
    // then use +8 to calcurate the vram address
    automatic logic signed [15:0] x = H_PixelCount - H_BackPorch + 8;
    automatic logic signed [15:0] y = V_PixelCount - V_BackPorch;
    logic active_area = (0 <= x && x < H_PixelValid + 8 && 0 <= y && y < V_PixelValid);

    if (!nRST) begin
      LCD_R <= 5'b00000;
      LCD_G <= 6'b000000;
      LCD_B <= 5'b00000;
    end else if (active_area) begin
      // get char code
      if (-2 <= x && x < H_PixelValid -2 + 8 && 0 <= y && y < V_PixelValid && (x+2) % 8 == 0) begin
        v_adb <= (x + 2) / 8 + (y / 16) * 60;
      end else if (-1 <= x && x < H_PixelValid -1 + 8 && 0 <= y && y < V_PixelValid && (x+1) % 8 == 0) begin
        char <= v_dout;
      end

      // draw the char
      // if (0 <= x && x < H_PixelValid && 0 <= y && y < V_PixelValid) begin
      if (char >= 0 && char <= 127) begin
        if (font[char][y%16][7-x%8] == 1'b1) begin
          LCD_R <= 5'b00000;  // green, foreground
          LCD_G <= 6'b111111;
          LCD_B <= 5'b00000;
        end else begin
          LCD_R <= 5'b00000;  // black, background
          LCD_G <= 6'b000000;
          LCD_B <= 5'b00000;
        end
      end else begin
        LCD_R <= 5'b11111;  // red (char is not defined)
        LCD_G <= 6'b000000;
        LCD_B <= 5'b00000;
      end
      // end else begin
      //   LCD_R <= 5'b00000;  // cyan (light blue)
      //   LCD_G <= 6'b111111;
      //   LCD_B <= 5'b11111;
      // end
    end else begin
      LCD_R <= 5'b11111;  // yellow
      LCD_G <= 6'b111111;
      LCD_B <= 5'b00000;
    end
  end

endmodule
