542: begin adb <= operands[15:0] + 8'h00 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
544: begin v_ada <= 544; v_din <= to_hexchar(dout[7:4]); end
545: begin v_ada <= 545; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h01 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
546: begin v_ada <= 546; v_din <= to_hexchar(dout[7:4]); end
547: begin v_ada <= 547; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h02 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
548: begin v_ada <= 548; v_din <= to_hexchar(dout[7:4]); end
549: begin v_ada <= 549; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h03 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
550: begin v_ada <= 550; v_din <= to_hexchar(dout[7:4]); end
551: begin v_ada <= 551; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h04 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
553: begin v_ada <= 553; v_din <= to_hexchar(dout[7:4]); end
554: begin v_ada <= 554; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h05 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
555: begin v_ada <= 555; v_din <= to_hexchar(dout[7:4]); end
556: begin v_ada <= 556; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h06 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
557: begin v_ada <= 557; v_din <= to_hexchar(dout[7:4]); end
558: begin v_ada <= 558; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h07 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
559: begin v_ada <= 559; v_din <= to_hexchar(dout[7:4]); end
560: begin v_ada <= 560; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h08 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
563: begin v_ada <= 563; v_din <= to_hexchar(dout[7:4]); end
564: begin v_ada <= 564; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h09 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
565: begin v_ada <= 565; v_din <= to_hexchar(dout[7:4]); end
566: begin v_ada <= 566; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h0A & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
567: begin v_ada <= 567; v_din <= to_hexchar(dout[7:4]); end
568: begin v_ada <= 568; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h0B & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
569: begin v_ada <= 569; v_din <= to_hexchar(dout[7:4]); end
570: begin v_ada <= 570; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h0C & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
572: begin v_ada <= 572; v_din <= to_hexchar(dout[7:4]); end
573: begin v_ada <= 573; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h0D & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
574: begin v_ada <= 574; v_din <= to_hexchar(dout[7:4]); end
575: begin v_ada <= 575; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h0E & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
576: begin v_ada <= 576; v_din <= to_hexchar(dout[7:4]); end
577: begin v_ada <= 577; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h0F & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z00; end
578: begin v_ada <= 578; v_din <= to_hexchar(dout[7:4]); end
579: begin v_ada <= 579; v_din <= to_hexchar(dout[3:0]); end
