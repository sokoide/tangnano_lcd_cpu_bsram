662: begin adb <= operands[15:0] + 8'h20 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
664: begin v_ada <= 664; v_din <= to_hexchar(dout[7:4]); end
665: begin v_ada <= 665; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h21 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
666: begin v_ada <= 666; v_din <= to_hexchar(dout[7:4]); end
667: begin v_ada <= 667; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h22 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
668: begin v_ada <= 668; v_din <= to_hexchar(dout[7:4]); end
669: begin v_ada <= 669; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h23 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
670: begin v_ada <= 670; v_din <= to_hexchar(dout[7:4]); end
671: begin v_ada <= 671; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h24 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
673: begin v_ada <= 673; v_din <= to_hexchar(dout[7:4]); end
674: begin v_ada <= 674; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h25 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
675: begin v_ada <= 675; v_din <= to_hexchar(dout[7:4]); end
676: begin v_ada <= 676; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h26 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
677: begin v_ada <= 677; v_din <= to_hexchar(dout[7:4]); end
678: begin v_ada <= 678; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h27 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
679: begin v_ada <= 679; v_din <= to_hexchar(dout[7:4]); end
680: begin v_ada <= 680; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h28 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
683: begin v_ada <= 683; v_din <= to_hexchar(dout[7:4]); end
684: begin v_ada <= 684; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h29 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
685: begin v_ada <= 685; v_din <= to_hexchar(dout[7:4]); end
686: begin v_ada <= 686; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h2A & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
687: begin v_ada <= 687; v_din <= to_hexchar(dout[7:4]); end
688: begin v_ada <= 688; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h2B & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
689: begin v_ada <= 689; v_din <= to_hexchar(dout[7:4]); end
690: begin v_ada <= 690; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h2C & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
692: begin v_ada <= 692; v_din <= to_hexchar(dout[7:4]); end
693: begin v_ada <= 693; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h2D & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
694: begin v_ada <= 694; v_din <= to_hexchar(dout[7:4]); end
695: begin v_ada <= 695; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h2E & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
696: begin v_ada <= 696; v_din <= to_hexchar(dout[7:4]); end
697: begin v_ada <= 697; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h2F & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
698: begin v_ada <= 698; v_din <= to_hexchar(dout[7:4]); end
699: begin v_ada <= 699; v_din <= to_hexchar(dout[3:0]); end
