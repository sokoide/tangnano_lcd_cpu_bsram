482: begin adb <= 8'h20; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
484: begin v_ada <= 484; v_din <= to_hexchar(dout[7:4]); end
485: begin v_ada <= 485; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h21; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
486: begin v_ada <= 486; v_din <= to_hexchar(dout[7:4]); end
487: begin v_ada <= 487; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h22; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
488: begin v_ada <= 488; v_din <= to_hexchar(dout[7:4]); end
489: begin v_ada <= 489; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h23; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
490: begin v_ada <= 490; v_din <= to_hexchar(dout[7:4]); end
491: begin v_ada <= 491; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h24; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
493: begin v_ada <= 493; v_din <= to_hexchar(dout[7:4]); end
494: begin v_ada <= 494; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h25; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
495: begin v_ada <= 495; v_din <= to_hexchar(dout[7:4]); end
496: begin v_ada <= 496; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h26; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
497: begin v_ada <= 497; v_din <= to_hexchar(dout[7:4]); end
498: begin v_ada <= 498; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h27; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
499: begin v_ada <= 499; v_din <= to_hexchar(dout[7:4]); end
500: begin v_ada <= 500; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h28; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
503: begin v_ada <= 503; v_din <= to_hexchar(dout[7:4]); end
504: begin v_ada <= 504; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h29; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
505: begin v_ada <= 505; v_din <= to_hexchar(dout[7:4]); end
506: begin v_ada <= 506; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h2A; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
507: begin v_ada <= 507; v_din <= to_hexchar(dout[7:4]); end
508: begin v_ada <= 508; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h2B; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
509: begin v_ada <= 509; v_din <= to_hexchar(dout[7:4]); end
510: begin v_ada <= 510; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h2C; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
512: begin v_ada <= 512; v_din <= to_hexchar(dout[7:4]); end
513: begin v_ada <= 513; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h2D; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
514: begin v_ada <= 514; v_din <= to_hexchar(dout[7:4]); end
515: begin v_ada <= 515; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h2E; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
516: begin v_ada <= 516; v_din <= to_hexchar(dout[7:4]); end
517: begin v_ada <= 517; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h2F; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z02; end
518: begin v_ada <= 518; v_din <= to_hexchar(dout[7:4]); end
519: begin v_ada <= 519; v_din <= to_hexchar(dout[3:0]); end
