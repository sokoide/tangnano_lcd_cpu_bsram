722: begin adb <= 8'h60; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
724: begin v_ada <= 724; v_din <= to_hexchar(dout[7:4]); end
725: begin v_ada <= 725; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h61; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
726: begin v_ada <= 726; v_din <= to_hexchar(dout[7:4]); end
727: begin v_ada <= 727; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h62; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
728: begin v_ada <= 728; v_din <= to_hexchar(dout[7:4]); end
729: begin v_ada <= 729; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h63; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
730: begin v_ada <= 730; v_din <= to_hexchar(dout[7:4]); end
731: begin v_ada <= 731; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h64; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
733: begin v_ada <= 733; v_din <= to_hexchar(dout[7:4]); end
734: begin v_ada <= 734; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h65; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
735: begin v_ada <= 735; v_din <= to_hexchar(dout[7:4]); end
736: begin v_ada <= 736; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h66; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
737: begin v_ada <= 737; v_din <= to_hexchar(dout[7:4]); end
738: begin v_ada <= 738; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h67; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
739: begin v_ada <= 739; v_din <= to_hexchar(dout[7:4]); end
740: begin v_ada <= 740; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h68; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
743: begin v_ada <= 743; v_din <= to_hexchar(dout[7:4]); end
744: begin v_ada <= 744; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h69; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
745: begin v_ada <= 745; v_din <= to_hexchar(dout[7:4]); end
746: begin v_ada <= 746; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h6A; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
747: begin v_ada <= 747; v_din <= to_hexchar(dout[7:4]); end
748: begin v_ada <= 748; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h6B; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
749: begin v_ada <= 749; v_din <= to_hexchar(dout[7:4]); end
750: begin v_ada <= 750; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h6C; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
752: begin v_ada <= 752; v_din <= to_hexchar(dout[7:4]); end
753: begin v_ada <= 753; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h6D; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
754: begin v_ada <= 754; v_din <= to_hexchar(dout[7:4]); end
755: begin v_ada <= 755; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h6E; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
756: begin v_ada <= 756; v_din <= to_hexchar(dout[7:4]); end
757: begin v_ada <= 757; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h6F; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z06; end
758: begin v_ada <= 758; v_din <= to_hexchar(dout[7:4]); end
759: begin v_ada <= 759; v_din <= to_hexchar(dout[3:0]); end
