logic [7:0] boot_program[256];

assign boot_program = '{
        0: 8'hA9,
        1: 8'h00,
        2: 8'h85,
        3: 8'h00,
        4: 8'hA9,
        5: 8'hE0,
        6: 8'h85,
        7: 8'h01,
        8: 8'hA9,
        9: 8'h00,
        10: 8'h8D,
        11: 8'h4E,
        12: 8'h02,
        13: 8'h8D,
        14: 8'h4F,
        15: 8'h02,
        16: 8'hFF,
        17: 8'h04,
        18: 8'h20,
        19: 8'h2F,
        20: 8'h02,
        21: 8'hEE,
        22: 8'h4E,
        23: 8'h02,
        24: 8'hD0,
        25: 8'h03,
        26: 8'hEE,
        27: 8'h4F,
        28: 8'h02,
        29: 8'hAD,
        30: 8'h4F,
        31: 8'h02,
        32: 8'hC9,
        33: 8'h04,
        34: 8'h90,
        35: 8'h08,
        36: 8'hA9,
        37: 8'h00,
        38: 8'h8D,
        39: 8'h4E,
        40: 8'h02,
        41: 8'h8D,
        42: 8'h4F,
        43: 8'h02,
        44: 8'h4C,
        45: 8'h10,
        46: 8'h02,
        47: 8'hA0,
        48: 8'h00,
        49: 8'hB9,
        50: 8'h50,
        51: 8'h02,
        52: 8'hF0,
        53: 8'h17,
        54: 8'hAD,
        55: 8'h4E,
        56: 8'h02,
        57: 8'h18,
        58: 8'h69,
        59: 8'h00,
        60: 8'h85,
        61: 8'h00,
        62: 8'hAD,
        63: 8'h4F,
        64: 8'h02,
        65: 8'h69,
        66: 8'hE0,
        67: 8'h85,
        68: 8'h01,
        69: 8'hB9,
        70: 8'h50,
        71: 8'h02,
        72: 8'h91,
        73: 8'h00,
        74: 8'hC8,
        75: 8'hD0,
        76: 8'hE7,
        77: 8'h60,
        78: 8'h00,
        79: 8'h00,
        80: 8'h20,
        81: 8'h48,
        82: 8'h65,
        83: 8'h6C,
        84: 8'h6C,
        85: 8'h6F,
        86: 8'h2C,
        87: 8'h20,
        88: 8'h57,
        89: 8'h6F,
        90: 8'h72,
        91: 8'h6C,
        92: 8'h64,
        93: 8'h21,
        94: 8'h00,
        default: 8'hEA
    };
parameter logic [7:0] boot_program_length = 95;
