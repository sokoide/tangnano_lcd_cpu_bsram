logic [7:0] boot_program[256];

assign boot_program = '{
        0: 8'hA9,
        1: 8'h00,
        2: 8'h85,
        3: 8'h00,
        4: 8'hA9,
        5: 8'hE0,
        6: 8'h85,
        7: 8'h01,
        8: 8'hA9,
        9: 8'h00,
        10: 8'h8D,
        11: 8'h4B,
        12: 8'h02,
        13: 8'h8D,
        14: 8'h4C,
        15: 8'h02,
        16: 8'hFF,
        17: 8'h04,
        18: 8'h20,
        19: 8'h2F,
        20: 8'h02,
        21: 8'hEE,
        22: 8'h4B,
        23: 8'h02,
        24: 8'hD0,
        25: 8'h03,
        26: 8'hEE,
        27: 8'h4C,
        28: 8'h02,
        29: 8'hAD,
        30: 8'h4C,
        31: 8'h02,
        32: 8'hC9,
        33: 8'h04,
        34: 8'h90,
        35: 8'h08,
        36: 8'hA9,
        37: 8'h00,
        38: 8'h8D,
        39: 8'h4B,
        40: 8'h02,
        41: 8'h8D,
        42: 8'h4C,
        43: 8'h02,
        44: 8'h4C,
        45: 8'h10,
        46: 8'h02,
        47: 8'hA0,
        48: 8'h00,
        49: 8'hAD,
        50: 8'h4B,
        51: 8'h02,
        52: 8'h18,
        53: 8'h69,
        54: 8'h00,
        55: 8'h85,
        56: 8'h00,
        57: 8'hAD,
        58: 8'h4C,
        59: 8'h02,
        60: 8'h69,
        61: 8'hE0,
        62: 8'h85,
        63: 8'h01,
        64: 8'hB9,
        65: 8'h4D,
        66: 8'h02,
        67: 8'hF0,
        68: 8'h05,
        69: 8'h91,
        70: 8'h00,
        71: 8'hC8,
        72: 8'hD0,
        73: 8'hE7,
        74: 8'h60,
        75: 8'h00,
        76: 8'h00,
        77: 8'h20,
        78: 8'h48,
        79: 8'h65,
        80: 8'h6C,
        81: 8'h6C,
        82: 8'h6F,
        83: 8'h2C,
        84: 8'h20,
        85: 8'h57,
        86: 8'h6F,
        87: 8'h72,
        88: 8'h6C,
        89: 8'h64,
        90: 8'h21,
        91: 8'h00,
        default: 8'hEA
    };
parameter logic [7:0] boot_program_length = 92;
