// Registers)
show_info_rom[0] = '{ v_ada: 10'd0, v_din_t: 2, v_din: 8'h52, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[1] = '{ v_ada: 10'd1, v_din_t: 2, v_din: 8'h65, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[2] = '{ v_ada: 10'd2, v_din_t: 2, v_din: 8'h67, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[3] = '{ v_ada: 10'd3, v_din_t: 2, v_din: 8'h69, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[4] = '{ v_ada: 10'd4, v_din_t: 2, v_din: 8'h73, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[5] = '{ v_ada: 10'd5, v_din_t: 2, v_din: 8'h74, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[6] = '{ v_ada: 10'd6, v_din_t: 2, v_din: 8'h65, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[7] = '{ v_ada: 10'd7, v_din_t: 2, v_din: 8'h72, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[8] = '{ v_ada: 10'd8, v_din_t: 2, v_din: 8'h73, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[9] = '{ v_ada: 10'd9, v_din_t: 2, v_din: 8'h29, diff: 8'h00, vram_write: 1, mem_read: 0};
// A :0x
show_info_rom[10] = '{ v_ada: 10'd60, v_din_t: 2, v_din: 8'h41, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[11] = '{ v_ada: 10'd61, v_din_t: 2, v_din: 8'h20, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[12] = '{ v_ada: 10'd62, v_din_t: 2, v_din: 8'h3A, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[13] = '{ v_ada: 10'd63, v_din_t: 2, v_din: 8'h30, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[14] = '{ v_ada: 10'd64, v_din_t: 2, v_din: 8'h78, diff: 8'h00, vram_write: 1, mem_read: 0};
// X :0x
show_info_rom[15] = '{ v_ada: 10'd120, v_din_t: 2, v_din: 8'h58, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[16] = '{ v_ada: 10'd121, v_din_t: 2, v_din: 8'h20, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[17] = '{ v_ada: 10'd122, v_din_t: 2, v_din: 8'h3A, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[18] = '{ v_ada: 10'd123, v_din_t: 2, v_din: 8'h30, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[19] = '{ v_ada: 10'd124, v_din_t: 2, v_din: 8'h78, diff: 8'h00, vram_write: 1, mem_read: 0};
// Y :0x
show_info_rom[20] = '{ v_ada: 10'd180, v_din_t: 2, v_din: 8'h59, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[21] = '{ v_ada: 10'd181, v_din_t: 2, v_din: 8'h20, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[22] = '{ v_ada: 10'd182, v_din_t: 2, v_din: 8'h3A, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[23] = '{ v_ada: 10'd183, v_din_t: 2, v_din: 8'h30, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[24] = '{ v_ada: 10'd184, v_din_t: 2, v_din: 8'h78, diff: 8'h00, vram_write: 1, mem_read: 0};
// PC:0x
show_info_rom[25] = '{ v_ada: 10'd240, v_din_t: 2, v_din: 8'h50, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[26] = '{ v_ada: 10'd241, v_din_t: 2, v_din: 8'h43, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[27] = '{ v_ada: 10'd242, v_din_t: 2, v_din: 8'h3A, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[28] = '{ v_ada: 10'd243, v_din_t: 2, v_din: 8'h30, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[29] = '{ v_ada: 10'd244, v_din_t: 2, v_din: 8'h78, diff: 8'h00, vram_write: 1, mem_read: 0};
// SP:0x
show_info_rom[30] = '{ v_ada: 10'd300, v_din_t: 2, v_din: 8'h53, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[31] = '{ v_ada: 10'd301, v_din_t: 2, v_din: 8'h50, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[32] = '{ v_ada: 10'd302, v_din_t: 2, v_din: 8'h3A, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[33] = '{ v_ada: 10'd303, v_din_t: 2, v_din: 8'h30, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[34] = '{ v_ada: 10'd304, v_din_t: 2, v_din: 8'h78, diff: 8'h00, vram_write: 1, mem_read: 0};
// Address 0x
show_info_rom[35] = '{ v_ada: 10'd480, v_din_t: 2, v_din: 8'h41, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[36] = '{ v_ada: 10'd481, v_din_t: 2, v_din: 8'h64, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[37] = '{ v_ada: 10'd482, v_din_t: 2, v_din: 8'h64, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[38] = '{ v_ada: 10'd483, v_din_t: 2, v_din: 8'h72, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[39] = '{ v_ada: 10'd484, v_din_t: 2, v_din: 8'h65, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[40] = '{ v_ada: 10'd485, v_din_t: 2, v_din: 8'h73, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[41] = '{ v_ada: 10'd486, v_din_t: 2, v_din: 8'h73, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[42] = '{ v_ada: 10'd487, v_din_t: 2, v_din: 8'h20, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[43] = '{ v_ada: 10'd488, v_din_t: 2, v_din: 8'h30, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[44] = '{ v_ada: 10'd489, v_din_t: 2, v_din: 8'h78, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[45] = '{ v_ada: 10'd490, v_din_t: 8, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[46] = '{ v_ada: 10'd491, v_din_t: 8, v_din: 8'h01, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[47] = '{ v_ada: 10'd492, v_din_t: 8, v_din: 8'h02, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[48] = '{ v_ada: 10'd493, v_din_t: 8, v_din: 8'h03, diff: 8'h00, vram_write: 1, mem_read: 0};
// -
show_info_rom[49] = '{ v_ada: 10'd494, v_din_t: 2, v_din: 8'h2D, diff: 8'h00, vram_write: 1, mem_read: 0};
// Memory dump
show_info_rom[50] = '{ v_ada: 10'd0, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 0, mem_read: 1};
show_info_rom[52] = '{ v_ada: 10'd544, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[53] = '{ v_ada: 10'd545, v_din_t: 1, v_din: 8'h00, diff: 8'h01, vram_write: 1, mem_read: 1};
show_info_rom[54] = '{ v_ada: 10'd546, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[55] = '{ v_ada: 10'd547, v_din_t: 1, v_din: 8'h00, diff: 8'h02, vram_write: 1, mem_read: 1};
show_info_rom[56] = '{ v_ada: 10'd548, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[57] = '{ v_ada: 10'd549, v_din_t: 1, v_din: 8'h00, diff: 8'h03, vram_write: 1, mem_read: 1};
show_info_rom[58] = '{ v_ada: 10'd550, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[59] = '{ v_ada: 10'd551, v_din_t: 1, v_din: 8'h00, diff: 8'h04, vram_write: 1, mem_read: 1};
show_info_rom[60] = '{ v_ada: 10'd553, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[61] = '{ v_ada: 10'd554, v_din_t: 1, v_din: 8'h00, diff: 8'h05, vram_write: 1, mem_read: 1};
show_info_rom[62] = '{ v_ada: 10'd555, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[63] = '{ v_ada: 10'd556, v_din_t: 1, v_din: 8'h00, diff: 8'h06, vram_write: 1, mem_read: 1};
show_info_rom[64] = '{ v_ada: 10'd557, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[65] = '{ v_ada: 10'd558, v_din_t: 1, v_din: 8'h00, diff: 8'h07, vram_write: 1, mem_read: 1};
show_info_rom[66] = '{ v_ada: 10'd559, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[67] = '{ v_ada: 10'd560, v_din_t: 1, v_din: 8'h00, diff: 8'h08, vram_write: 1, mem_read: 1};
show_info_rom[68] = '{ v_ada: 10'd563, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[69] = '{ v_ada: 10'd564, v_din_t: 1, v_din: 8'h00, diff: 8'h09, vram_write: 1, mem_read: 1};
show_info_rom[70] = '{ v_ada: 10'd565, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[71] = '{ v_ada: 10'd566, v_din_t: 1, v_din: 8'h00, diff: 8'h0A, vram_write: 1, mem_read: 1};
show_info_rom[72] = '{ v_ada: 10'd567, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[73] = '{ v_ada: 10'd568, v_din_t: 1, v_din: 8'h00, diff: 8'h0B, vram_write: 1, mem_read: 1};
show_info_rom[74] = '{ v_ada: 10'd569, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[75] = '{ v_ada: 10'd570, v_din_t: 1, v_din: 8'h00, diff: 8'h0C, vram_write: 1, mem_read: 1};
show_info_rom[76] = '{ v_ada: 10'd572, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[77] = '{ v_ada: 10'd573, v_din_t: 1, v_din: 8'h00, diff: 8'h0D, vram_write: 1, mem_read: 1};
show_info_rom[78] = '{ v_ada: 10'd574, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[79] = '{ v_ada: 10'd575, v_din_t: 1, v_din: 8'h00, diff: 8'h0E, vram_write: 1, mem_read: 1};
show_info_rom[80] = '{ v_ada: 10'd576, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[81] = '{ v_ada: 10'd577, v_din_t: 1, v_din: 8'h00, diff: 8'h0F, vram_write: 1, mem_read: 1};
show_info_rom[82] = '{ v_ada: 10'd578, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[83] = '{ v_ada: 10'd579, v_din_t: 1, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[84] = '{ v_ada: 10'd0, v_din_t: 0, v_din: 8'h00, diff: 8'h10, vram_write: 0, mem_read: 1};
show_info_rom[86] = '{ v_ada: 10'd604, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[87] = '{ v_ada: 10'd605, v_din_t: 1, v_din: 8'h00, diff: 8'h11, vram_write: 1, mem_read: 1};
show_info_rom[88] = '{ v_ada: 10'd606, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[89] = '{ v_ada: 10'd607, v_din_t: 1, v_din: 8'h00, diff: 8'h12, vram_write: 1, mem_read: 1};
show_info_rom[90] = '{ v_ada: 10'd608, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[91] = '{ v_ada: 10'd609, v_din_t: 1, v_din: 8'h00, diff: 8'h13, vram_write: 1, mem_read: 1};
show_info_rom[92] = '{ v_ada: 10'd610, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[93] = '{ v_ada: 10'd611, v_din_t: 1, v_din: 8'h00, diff: 8'h14, vram_write: 1, mem_read: 1};
show_info_rom[94] = '{ v_ada: 10'd613, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[95] = '{ v_ada: 10'd614, v_din_t: 1, v_din: 8'h00, diff: 8'h15, vram_write: 1, mem_read: 1};
show_info_rom[96] = '{ v_ada: 10'd615, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[97] = '{ v_ada: 10'd616, v_din_t: 1, v_din: 8'h00, diff: 8'h16, vram_write: 1, mem_read: 1};
show_info_rom[98] = '{ v_ada: 10'd617, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[99] = '{ v_ada: 10'd618, v_din_t: 1, v_din: 8'h00, diff: 8'h17, vram_write: 1, mem_read: 1};
show_info_rom[100] = '{ v_ada: 10'd619, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[101] = '{ v_ada: 10'd620, v_din_t: 1, v_din: 8'h00, diff: 8'h18, vram_write: 1, mem_read: 1};
show_info_rom[102] = '{ v_ada: 10'd623, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[103] = '{ v_ada: 10'd624, v_din_t: 1, v_din: 8'h00, diff: 8'h19, vram_write: 1, mem_read: 1};
show_info_rom[104] = '{ v_ada: 10'd625, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[105] = '{ v_ada: 10'd626, v_din_t: 1, v_din: 8'h00, diff: 8'h1A, vram_write: 1, mem_read: 1};
show_info_rom[106] = '{ v_ada: 10'd627, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[107] = '{ v_ada: 10'd628, v_din_t: 1, v_din: 8'h00, diff: 8'h1B, vram_write: 1, mem_read: 1};
show_info_rom[108] = '{ v_ada: 10'd629, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[109] = '{ v_ada: 10'd630, v_din_t: 1, v_din: 8'h00, diff: 8'h1C, vram_write: 1, mem_read: 1};
show_info_rom[110] = '{ v_ada: 10'd632, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[111] = '{ v_ada: 10'd633, v_din_t: 1, v_din: 8'h00, diff: 8'h1D, vram_write: 1, mem_read: 1};
show_info_rom[112] = '{ v_ada: 10'd634, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[113] = '{ v_ada: 10'd635, v_din_t: 1, v_din: 8'h00, diff: 8'h1E, vram_write: 1, mem_read: 1};
show_info_rom[114] = '{ v_ada: 10'd636, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[115] = '{ v_ada: 10'd637, v_din_t: 1, v_din: 8'h00, diff: 8'h1F, vram_write: 1, mem_read: 1};
show_info_rom[116] = '{ v_ada: 10'd638, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[117] = '{ v_ada: 10'd639, v_din_t: 1, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[118] = '{ v_ada: 10'd0, v_din_t: 0, v_din: 8'h00, diff: 8'h20, vram_write: 0, mem_read: 1};
show_info_rom[120] = '{ v_ada: 10'd664, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[121] = '{ v_ada: 10'd665, v_din_t: 1, v_din: 8'h00, diff: 8'h21, vram_write: 1, mem_read: 1};
show_info_rom[122] = '{ v_ada: 10'd666, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[123] = '{ v_ada: 10'd667, v_din_t: 1, v_din: 8'h00, diff: 8'h22, vram_write: 1, mem_read: 1};
show_info_rom[124] = '{ v_ada: 10'd668, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[125] = '{ v_ada: 10'd669, v_din_t: 1, v_din: 8'h00, diff: 8'h23, vram_write: 1, mem_read: 1};
show_info_rom[126] = '{ v_ada: 10'd670, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[127] = '{ v_ada: 10'd671, v_din_t: 1, v_din: 8'h00, diff: 8'h24, vram_write: 1, mem_read: 1};
show_info_rom[128] = '{ v_ada: 10'd673, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[129] = '{ v_ada: 10'd674, v_din_t: 1, v_din: 8'h00, diff: 8'h25, vram_write: 1, mem_read: 1};
show_info_rom[130] = '{ v_ada: 10'd675, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[131] = '{ v_ada: 10'd676, v_din_t: 1, v_din: 8'h00, diff: 8'h26, vram_write: 1, mem_read: 1};
show_info_rom[132] = '{ v_ada: 10'd677, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[133] = '{ v_ada: 10'd678, v_din_t: 1, v_din: 8'h00, diff: 8'h27, vram_write: 1, mem_read: 1};
show_info_rom[134] = '{ v_ada: 10'd679, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[135] = '{ v_ada: 10'd680, v_din_t: 1, v_din: 8'h00, diff: 8'h28, vram_write: 1, mem_read: 1};
show_info_rom[136] = '{ v_ada: 10'd683, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[137] = '{ v_ada: 10'd684, v_din_t: 1, v_din: 8'h00, diff: 8'h29, vram_write: 1, mem_read: 1};
show_info_rom[138] = '{ v_ada: 10'd685, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[139] = '{ v_ada: 10'd686, v_din_t: 1, v_din: 8'h00, diff: 8'h2A, vram_write: 1, mem_read: 1};
show_info_rom[140] = '{ v_ada: 10'd687, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[141] = '{ v_ada: 10'd688, v_din_t: 1, v_din: 8'h00, diff: 8'h2B, vram_write: 1, mem_read: 1};
show_info_rom[142] = '{ v_ada: 10'd689, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[143] = '{ v_ada: 10'd690, v_din_t: 1, v_din: 8'h00, diff: 8'h2C, vram_write: 1, mem_read: 1};
show_info_rom[144] = '{ v_ada: 10'd692, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[145] = '{ v_ada: 10'd693, v_din_t: 1, v_din: 8'h00, diff: 8'h2D, vram_write: 1, mem_read: 1};
show_info_rom[146] = '{ v_ada: 10'd694, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[147] = '{ v_ada: 10'd695, v_din_t: 1, v_din: 8'h00, diff: 8'h2E, vram_write: 1, mem_read: 1};
show_info_rom[148] = '{ v_ada: 10'd696, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[149] = '{ v_ada: 10'd697, v_din_t: 1, v_din: 8'h00, diff: 8'h2F, vram_write: 1, mem_read: 1};
show_info_rom[150] = '{ v_ada: 10'd698, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[151] = '{ v_ada: 10'd699, v_din_t: 1, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[152] = '{ v_ada: 10'd0, v_din_t: 0, v_din: 8'h00, diff: 8'h30, vram_write: 0, mem_read: 1};
show_info_rom[154] = '{ v_ada: 10'd724, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[155] = '{ v_ada: 10'd725, v_din_t: 1, v_din: 8'h00, diff: 8'h31, vram_write: 1, mem_read: 1};
show_info_rom[156] = '{ v_ada: 10'd726, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[157] = '{ v_ada: 10'd727, v_din_t: 1, v_din: 8'h00, diff: 8'h32, vram_write: 1, mem_read: 1};
show_info_rom[158] = '{ v_ada: 10'd728, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[159] = '{ v_ada: 10'd729, v_din_t: 1, v_din: 8'h00, diff: 8'h33, vram_write: 1, mem_read: 1};
show_info_rom[160] = '{ v_ada: 10'd730, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[161] = '{ v_ada: 10'd731, v_din_t: 1, v_din: 8'h00, diff: 8'h34, vram_write: 1, mem_read: 1};
show_info_rom[162] = '{ v_ada: 10'd733, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[163] = '{ v_ada: 10'd734, v_din_t: 1, v_din: 8'h00, diff: 8'h35, vram_write: 1, mem_read: 1};
show_info_rom[164] = '{ v_ada: 10'd735, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[165] = '{ v_ada: 10'd736, v_din_t: 1, v_din: 8'h00, diff: 8'h36, vram_write: 1, mem_read: 1};
show_info_rom[166] = '{ v_ada: 10'd737, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[167] = '{ v_ada: 10'd738, v_din_t: 1, v_din: 8'h00, diff: 8'h37, vram_write: 1, mem_read: 1};
show_info_rom[168] = '{ v_ada: 10'd739, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[169] = '{ v_ada: 10'd740, v_din_t: 1, v_din: 8'h00, diff: 8'h38, vram_write: 1, mem_read: 1};
show_info_rom[170] = '{ v_ada: 10'd743, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[171] = '{ v_ada: 10'd744, v_din_t: 1, v_din: 8'h00, diff: 8'h39, vram_write: 1, mem_read: 1};
show_info_rom[172] = '{ v_ada: 10'd745, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[173] = '{ v_ada: 10'd746, v_din_t: 1, v_din: 8'h00, diff: 8'h3A, vram_write: 1, mem_read: 1};
show_info_rom[174] = '{ v_ada: 10'd747, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[175] = '{ v_ada: 10'd748, v_din_t: 1, v_din: 8'h00, diff: 8'h3B, vram_write: 1, mem_read: 1};
show_info_rom[176] = '{ v_ada: 10'd749, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[177] = '{ v_ada: 10'd750, v_din_t: 1, v_din: 8'h00, diff: 8'h3C, vram_write: 1, mem_read: 1};
show_info_rom[178] = '{ v_ada: 10'd752, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[179] = '{ v_ada: 10'd753, v_din_t: 1, v_din: 8'h00, diff: 8'h3D, vram_write: 1, mem_read: 1};
show_info_rom[180] = '{ v_ada: 10'd754, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[181] = '{ v_ada: 10'd755, v_din_t: 1, v_din: 8'h00, diff: 8'h3E, vram_write: 1, mem_read: 1};
show_info_rom[182] = '{ v_ada: 10'd756, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[183] = '{ v_ada: 10'd757, v_din_t: 1, v_din: 8'h00, diff: 8'h3F, vram_write: 1, mem_read: 1};
show_info_rom[184] = '{ v_ada: 10'd758, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[185] = '{ v_ada: 10'd759, v_din_t: 1, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[186] = '{ v_ada: 10'd0, v_din_t: 0, v_din: 8'h00, diff: 8'h40, vram_write: 0, mem_read: 1};
show_info_rom[188] = '{ v_ada: 10'd784, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[189] = '{ v_ada: 10'd785, v_din_t: 1, v_din: 8'h00, diff: 8'h41, vram_write: 1, mem_read: 1};
show_info_rom[190] = '{ v_ada: 10'd786, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[191] = '{ v_ada: 10'd787, v_din_t: 1, v_din: 8'h00, diff: 8'h42, vram_write: 1, mem_read: 1};
show_info_rom[192] = '{ v_ada: 10'd788, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[193] = '{ v_ada: 10'd789, v_din_t: 1, v_din: 8'h00, diff: 8'h43, vram_write: 1, mem_read: 1};
show_info_rom[194] = '{ v_ada: 10'd790, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[195] = '{ v_ada: 10'd791, v_din_t: 1, v_din: 8'h00, diff: 8'h44, vram_write: 1, mem_read: 1};
show_info_rom[196] = '{ v_ada: 10'd793, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[197] = '{ v_ada: 10'd794, v_din_t: 1, v_din: 8'h00, diff: 8'h45, vram_write: 1, mem_read: 1};
show_info_rom[198] = '{ v_ada: 10'd795, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[199] = '{ v_ada: 10'd796, v_din_t: 1, v_din: 8'h00, diff: 8'h46, vram_write: 1, mem_read: 1};
show_info_rom[200] = '{ v_ada: 10'd797, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[201] = '{ v_ada: 10'd798, v_din_t: 1, v_din: 8'h00, diff: 8'h47, vram_write: 1, mem_read: 1};
show_info_rom[202] = '{ v_ada: 10'd799, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[203] = '{ v_ada: 10'd800, v_din_t: 1, v_din: 8'h00, diff: 8'h48, vram_write: 1, mem_read: 1};
show_info_rom[204] = '{ v_ada: 10'd803, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[205] = '{ v_ada: 10'd804, v_din_t: 1, v_din: 8'h00, diff: 8'h49, vram_write: 1, mem_read: 1};
show_info_rom[206] = '{ v_ada: 10'd805, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[207] = '{ v_ada: 10'd806, v_din_t: 1, v_din: 8'h00, diff: 8'h4A, vram_write: 1, mem_read: 1};
show_info_rom[208] = '{ v_ada: 10'd807, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[209] = '{ v_ada: 10'd808, v_din_t: 1, v_din: 8'h00, diff: 8'h4B, vram_write: 1, mem_read: 1};
show_info_rom[210] = '{ v_ada: 10'd809, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[211] = '{ v_ada: 10'd810, v_din_t: 1, v_din: 8'h00, diff: 8'h4C, vram_write: 1, mem_read: 1};
show_info_rom[212] = '{ v_ada: 10'd812, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[213] = '{ v_ada: 10'd813, v_din_t: 1, v_din: 8'h00, diff: 8'h4D, vram_write: 1, mem_read: 1};
show_info_rom[214] = '{ v_ada: 10'd814, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[215] = '{ v_ada: 10'd815, v_din_t: 1, v_din: 8'h00, diff: 8'h4E, vram_write: 1, mem_read: 1};
show_info_rom[216] = '{ v_ada: 10'd816, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[217] = '{ v_ada: 10'd817, v_din_t: 1, v_din: 8'h00, diff: 8'h4F, vram_write: 1, mem_read: 1};
show_info_rom[218] = '{ v_ada: 10'd818, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[219] = '{ v_ada: 10'd819, v_din_t: 1, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[220] = '{ v_ada: 10'd0, v_din_t: 0, v_din: 8'h00, diff: 8'h50, vram_write: 0, mem_read: 1};
show_info_rom[222] = '{ v_ada: 10'd844, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[223] = '{ v_ada: 10'd845, v_din_t: 1, v_din: 8'h00, diff: 8'h51, vram_write: 1, mem_read: 1};
show_info_rom[224] = '{ v_ada: 10'd846, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[225] = '{ v_ada: 10'd847, v_din_t: 1, v_din: 8'h00, diff: 8'h52, vram_write: 1, mem_read: 1};
show_info_rom[226] = '{ v_ada: 10'd848, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[227] = '{ v_ada: 10'd849, v_din_t: 1, v_din: 8'h00, diff: 8'h53, vram_write: 1, mem_read: 1};
show_info_rom[228] = '{ v_ada: 10'd850, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[229] = '{ v_ada: 10'd851, v_din_t: 1, v_din: 8'h00, diff: 8'h54, vram_write: 1, mem_read: 1};
show_info_rom[230] = '{ v_ada: 10'd853, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[231] = '{ v_ada: 10'd854, v_din_t: 1, v_din: 8'h00, diff: 8'h55, vram_write: 1, mem_read: 1};
show_info_rom[232] = '{ v_ada: 10'd855, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[233] = '{ v_ada: 10'd856, v_din_t: 1, v_din: 8'h00, diff: 8'h56, vram_write: 1, mem_read: 1};
show_info_rom[234] = '{ v_ada: 10'd857, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[235] = '{ v_ada: 10'd858, v_din_t: 1, v_din: 8'h00, diff: 8'h57, vram_write: 1, mem_read: 1};
show_info_rom[236] = '{ v_ada: 10'd859, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[237] = '{ v_ada: 10'd860, v_din_t: 1, v_din: 8'h00, diff: 8'h58, vram_write: 1, mem_read: 1};
show_info_rom[238] = '{ v_ada: 10'd863, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[239] = '{ v_ada: 10'd864, v_din_t: 1, v_din: 8'h00, diff: 8'h59, vram_write: 1, mem_read: 1};
show_info_rom[240] = '{ v_ada: 10'd865, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[241] = '{ v_ada: 10'd866, v_din_t: 1, v_din: 8'h00, diff: 8'h5A, vram_write: 1, mem_read: 1};
show_info_rom[242] = '{ v_ada: 10'd867, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[243] = '{ v_ada: 10'd868, v_din_t: 1, v_din: 8'h00, diff: 8'h5B, vram_write: 1, mem_read: 1};
show_info_rom[244] = '{ v_ada: 10'd869, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[245] = '{ v_ada: 10'd870, v_din_t: 1, v_din: 8'h00, diff: 8'h5C, vram_write: 1, mem_read: 1};
show_info_rom[246] = '{ v_ada: 10'd872, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[247] = '{ v_ada: 10'd873, v_din_t: 1, v_din: 8'h00, diff: 8'h5D, vram_write: 1, mem_read: 1};
show_info_rom[248] = '{ v_ada: 10'd874, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[249] = '{ v_ada: 10'd875, v_din_t: 1, v_din: 8'h00, diff: 8'h5E, vram_write: 1, mem_read: 1};
show_info_rom[250] = '{ v_ada: 10'd876, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[251] = '{ v_ada: 10'd877, v_din_t: 1, v_din: 8'h00, diff: 8'h5F, vram_write: 1, mem_read: 1};
show_info_rom[252] = '{ v_ada: 10'd878, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[253] = '{ v_ada: 10'd879, v_din_t: 1, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[254] = '{ v_ada: 10'd0, v_din_t: 0, v_din: 8'h00, diff: 8'h60, vram_write: 0, mem_read: 1};
show_info_rom[256] = '{ v_ada: 10'd904, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[257] = '{ v_ada: 10'd905, v_din_t: 1, v_din: 8'h00, diff: 8'h61, vram_write: 1, mem_read: 1};
show_info_rom[258] = '{ v_ada: 10'd906, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[259] = '{ v_ada: 10'd907, v_din_t: 1, v_din: 8'h00, diff: 8'h62, vram_write: 1, mem_read: 1};
show_info_rom[260] = '{ v_ada: 10'd908, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[261] = '{ v_ada: 10'd909, v_din_t: 1, v_din: 8'h00, diff: 8'h63, vram_write: 1, mem_read: 1};
show_info_rom[262] = '{ v_ada: 10'd910, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[263] = '{ v_ada: 10'd911, v_din_t: 1, v_din: 8'h00, diff: 8'h64, vram_write: 1, mem_read: 1};
show_info_rom[264] = '{ v_ada: 10'd913, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[265] = '{ v_ada: 10'd914, v_din_t: 1, v_din: 8'h00, diff: 8'h65, vram_write: 1, mem_read: 1};
show_info_rom[266] = '{ v_ada: 10'd915, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[267] = '{ v_ada: 10'd916, v_din_t: 1, v_din: 8'h00, diff: 8'h66, vram_write: 1, mem_read: 1};
show_info_rom[268] = '{ v_ada: 10'd917, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[269] = '{ v_ada: 10'd918, v_din_t: 1, v_din: 8'h00, diff: 8'h67, vram_write: 1, mem_read: 1};
show_info_rom[270] = '{ v_ada: 10'd919, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[271] = '{ v_ada: 10'd920, v_din_t: 1, v_din: 8'h00, diff: 8'h68, vram_write: 1, mem_read: 1};
show_info_rom[272] = '{ v_ada: 10'd923, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[273] = '{ v_ada: 10'd924, v_din_t: 1, v_din: 8'h00, diff: 8'h69, vram_write: 1, mem_read: 1};
show_info_rom[274] = '{ v_ada: 10'd925, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[275] = '{ v_ada: 10'd926, v_din_t: 1, v_din: 8'h00, diff: 8'h6A, vram_write: 1, mem_read: 1};
show_info_rom[276] = '{ v_ada: 10'd927, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[277] = '{ v_ada: 10'd928, v_din_t: 1, v_din: 8'h00, diff: 8'h6B, vram_write: 1, mem_read: 1};
show_info_rom[278] = '{ v_ada: 10'd929, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[279] = '{ v_ada: 10'd930, v_din_t: 1, v_din: 8'h00, diff: 8'h6C, vram_write: 1, mem_read: 1};
show_info_rom[280] = '{ v_ada: 10'd932, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[281] = '{ v_ada: 10'd933, v_din_t: 1, v_din: 8'h00, diff: 8'h6D, vram_write: 1, mem_read: 1};
show_info_rom[282] = '{ v_ada: 10'd934, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[283] = '{ v_ada: 10'd935, v_din_t: 1, v_din: 8'h00, diff: 8'h6E, vram_write: 1, mem_read: 1};
show_info_rom[284] = '{ v_ada: 10'd936, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[285] = '{ v_ada: 10'd937, v_din_t: 1, v_din: 8'h00, diff: 8'h6F, vram_write: 1, mem_read: 1};
show_info_rom[286] = '{ v_ada: 10'd938, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[287] = '{ v_ada: 10'd939, v_din_t: 1, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[288] = '{ v_ada: 10'd0, v_din_t: 0, v_din: 8'h00, diff: 8'h70, vram_write: 0, mem_read: 1};
show_info_rom[290] = '{ v_ada: 10'd964, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[291] = '{ v_ada: 10'd965, v_din_t: 1, v_din: 8'h00, diff: 8'h71, vram_write: 1, mem_read: 1};
show_info_rom[292] = '{ v_ada: 10'd966, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[293] = '{ v_ada: 10'd967, v_din_t: 1, v_din: 8'h00, diff: 8'h72, vram_write: 1, mem_read: 1};
show_info_rom[294] = '{ v_ada: 10'd968, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[295] = '{ v_ada: 10'd969, v_din_t: 1, v_din: 8'h00, diff: 8'h73, vram_write: 1, mem_read: 1};
show_info_rom[296] = '{ v_ada: 10'd970, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[297] = '{ v_ada: 10'd971, v_din_t: 1, v_din: 8'h00, diff: 8'h74, vram_write: 1, mem_read: 1};
show_info_rom[298] = '{ v_ada: 10'd973, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[299] = '{ v_ada: 10'd974, v_din_t: 1, v_din: 8'h00, diff: 8'h75, vram_write: 1, mem_read: 1};
show_info_rom[300] = '{ v_ada: 10'd975, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[301] = '{ v_ada: 10'd976, v_din_t: 1, v_din: 8'h00, diff: 8'h76, vram_write: 1, mem_read: 1};
show_info_rom[302] = '{ v_ada: 10'd977, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[303] = '{ v_ada: 10'd978, v_din_t: 1, v_din: 8'h00, diff: 8'h77, vram_write: 1, mem_read: 1};
show_info_rom[304] = '{ v_ada: 10'd979, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[305] = '{ v_ada: 10'd980, v_din_t: 1, v_din: 8'h00, diff: 8'h78, vram_write: 1, mem_read: 1};
show_info_rom[306] = '{ v_ada: 10'd983, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[307] = '{ v_ada: 10'd984, v_din_t: 1, v_din: 8'h00, diff: 8'h79, vram_write: 1, mem_read: 1};
show_info_rom[308] = '{ v_ada: 10'd985, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[309] = '{ v_ada: 10'd986, v_din_t: 1, v_din: 8'h00, diff: 8'h7A, vram_write: 1, mem_read: 1};
show_info_rom[310] = '{ v_ada: 10'd987, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[311] = '{ v_ada: 10'd988, v_din_t: 1, v_din: 8'h00, diff: 8'h7B, vram_write: 1, mem_read: 1};
show_info_rom[312] = '{ v_ada: 10'd989, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[313] = '{ v_ada: 10'd990, v_din_t: 1, v_din: 8'h00, diff: 8'h7C, vram_write: 1, mem_read: 1};
show_info_rom[314] = '{ v_ada: 10'd992, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[315] = '{ v_ada: 10'd993, v_din_t: 1, v_din: 8'h00, diff: 8'h7D, vram_write: 1, mem_read: 1};
show_info_rom[316] = '{ v_ada: 10'd994, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[317] = '{ v_ada: 10'd995, v_din_t: 1, v_din: 8'h00, diff: 8'h7E, vram_write: 1, mem_read: 1};
show_info_rom[318] = '{ v_ada: 10'd996, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[319] = '{ v_ada: 10'd997, v_din_t: 1, v_din: 8'h00, diff: 8'h7F, vram_write: 1, mem_read: 1};
show_info_rom[320] = '{ v_ada: 10'd998, v_din_t: 0, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
show_info_rom[321] = '{ v_ada: 10'd999, v_din_t: 1, v_din: 8'h00, diff: 8'h00, vram_write: 1, mem_read: 0};
