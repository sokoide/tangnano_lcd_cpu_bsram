`include "consts.svh"

module cpu();


endmodule