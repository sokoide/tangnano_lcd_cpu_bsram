662: begin adb <= 8'h50; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
664: begin v_ada <= 664; v_din <= to_hexchar(dout[7:4]); end
665: begin v_ada <= 665; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h51; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
666: begin v_ada <= 666; v_din <= to_hexchar(dout[7:4]); end
667: begin v_ada <= 667; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h52; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
668: begin v_ada <= 668; v_din <= to_hexchar(dout[7:4]); end
669: begin v_ada <= 669; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h53; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
670: begin v_ada <= 670; v_din <= to_hexchar(dout[7:4]); end
671: begin v_ada <= 671; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h54; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
673: begin v_ada <= 673; v_din <= to_hexchar(dout[7:4]); end
674: begin v_ada <= 674; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h55; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
675: begin v_ada <= 675; v_din <= to_hexchar(dout[7:4]); end
676: begin v_ada <= 676; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h56; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
677: begin v_ada <= 677; v_din <= to_hexchar(dout[7:4]); end
678: begin v_ada <= 678; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h57; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
679: begin v_ada <= 679; v_din <= to_hexchar(dout[7:4]); end
680: begin v_ada <= 680; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h58; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
683: begin v_ada <= 683; v_din <= to_hexchar(dout[7:4]); end
684: begin v_ada <= 684; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h59; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
685: begin v_ada <= 685; v_din <= to_hexchar(dout[7:4]); end
686: begin v_ada <= 686; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h5A; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
687: begin v_ada <= 687; v_din <= to_hexchar(dout[7:4]); end
688: begin v_ada <= 688; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h5B; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
689: begin v_ada <= 689; v_din <= to_hexchar(dout[7:4]); end
690: begin v_ada <= 690; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h5C; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
692: begin v_ada <= 692; v_din <= to_hexchar(dout[7:4]); end
693: begin v_ada <= 693; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h5D; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
694: begin v_ada <= 694; v_din <= to_hexchar(dout[7:4]); end
695: begin v_ada <= 695; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h5E; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
696: begin v_ada <= 696; v_din <= to_hexchar(dout[7:4]); end
697: begin v_ada <= 697; v_din <= to_hexchar(dout[3:0]);  adb <= 8'h5F; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
698: begin v_ada <= 698; v_din <= to_hexchar(dout[7:4]); end
699: begin v_ada <= 699; v_din <= to_hexchar(dout[3:0]); end
