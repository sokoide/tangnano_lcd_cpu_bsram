842: begin adb <= operands[15:0] + 8'h50 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
844: begin v_ada <= 844; v_din <= to_hexchar(dout[7:4]); end
845: begin v_ada <= 845; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h51 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
846: begin v_ada <= 846; v_din <= to_hexchar(dout[7:4]); end
847: begin v_ada <= 847; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h52 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
848: begin v_ada <= 848; v_din <= to_hexchar(dout[7:4]); end
849: begin v_ada <= 849; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h53 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
850: begin v_ada <= 850; v_din <= to_hexchar(dout[7:4]); end
851: begin v_ada <= 851; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h54 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
853: begin v_ada <= 853; v_din <= to_hexchar(dout[7:4]); end
854: begin v_ada <= 854; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h55 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
855: begin v_ada <= 855; v_din <= to_hexchar(dout[7:4]); end
856: begin v_ada <= 856; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h56 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
857: begin v_ada <= 857; v_din <= to_hexchar(dout[7:4]); end
858: begin v_ada <= 858; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h57 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
859: begin v_ada <= 859; v_din <= to_hexchar(dout[7:4]); end
860: begin v_ada <= 860; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h58 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
863: begin v_ada <= 863; v_din <= to_hexchar(dout[7:4]); end
864: begin v_ada <= 864; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h59 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
865: begin v_ada <= 865; v_din <= to_hexchar(dout[7:4]); end
866: begin v_ada <= 866; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h5A & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
867: begin v_ada <= 867; v_din <= to_hexchar(dout[7:4]); end
868: begin v_ada <= 868; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h5B & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
869: begin v_ada <= 869; v_din <= to_hexchar(dout[7:4]); end
870: begin v_ada <= 870; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h5C & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
872: begin v_ada <= 872; v_din <= to_hexchar(dout[7:4]); end
873: begin v_ada <= 873; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h5D & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
874: begin v_ada <= 874; v_din <= to_hexchar(dout[7:4]); end
875: begin v_ada <= 875; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h5E & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
876: begin v_ada <= 876; v_din <= to_hexchar(dout[7:4]); end
877: begin v_ada <= 877; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h5F & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z05; end
878: begin v_ada <= 878; v_din <= to_hexchar(dout[7:4]); end
879: begin v_ada <= 879; v_din <= to_hexchar(dout[3:0]); end
