602: begin adb <= operands[15:0] + 8'h10 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
604: begin v_ada <= 604; v_din <= to_hexchar(dout[7:4]); end
605: begin v_ada <= 605; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h11 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
606: begin v_ada <= 606; v_din <= to_hexchar(dout[7:4]); end
607: begin v_ada <= 607; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h12 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
608: begin v_ada <= 608; v_din <= to_hexchar(dout[7:4]); end
609: begin v_ada <= 609; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h13 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
610: begin v_ada <= 610; v_din <= to_hexchar(dout[7:4]); end
611: begin v_ada <= 611; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h14 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
613: begin v_ada <= 613; v_din <= to_hexchar(dout[7:4]); end
614: begin v_ada <= 614; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h15 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
615: begin v_ada <= 615; v_din <= to_hexchar(dout[7:4]); end
616: begin v_ada <= 616; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h16 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
617: begin v_ada <= 617; v_din <= to_hexchar(dout[7:4]); end
618: begin v_ada <= 618; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h17 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
619: begin v_ada <= 619; v_din <= to_hexchar(dout[7:4]); end
620: begin v_ada <= 620; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h18 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
623: begin v_ada <= 623; v_din <= to_hexchar(dout[7:4]); end
624: begin v_ada <= 624; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h19 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
625: begin v_ada <= 625; v_din <= to_hexchar(dout[7:4]); end
626: begin v_ada <= 626; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h1A & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
627: begin v_ada <= 627; v_din <= to_hexchar(dout[7:4]); end
628: begin v_ada <= 628; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h1B & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
629: begin v_ada <= 629; v_din <= to_hexchar(dout[7:4]); end
630: begin v_ada <= 630; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h1C & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
632: begin v_ada <= 632; v_din <= to_hexchar(dout[7:4]); end
633: begin v_ada <= 633; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h1D & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
634: begin v_ada <= 634; v_din <= to_hexchar(dout[7:4]); end
635: begin v_ada <= 635; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h1E & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
636: begin v_ada <= 636; v_din <= to_hexchar(dout[7:4]); end
637: begin v_ada <= 637; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h1F & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z01; end
638: begin v_ada <= 638; v_din <= to_hexchar(dout[7:4]); end
639: begin v_ada <= 639; v_din <= to_hexchar(dout[3:0]); end
