module cpu();


endmodule