962: begin adb <= operands[15:0] + 8'h70 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
964: begin v_ada <= 964; v_din <= to_hexchar(dout[7:4]); end
965: begin v_ada <= 965; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h71 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
966: begin v_ada <= 966; v_din <= to_hexchar(dout[7:4]); end
967: begin v_ada <= 967; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h72 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
968: begin v_ada <= 968; v_din <= to_hexchar(dout[7:4]); end
969: begin v_ada <= 969; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h73 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
970: begin v_ada <= 970; v_din <= to_hexchar(dout[7:4]); end
971: begin v_ada <= 971; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h74 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
973: begin v_ada <= 973; v_din <= to_hexchar(dout[7:4]); end
974: begin v_ada <= 974; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h75 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
975: begin v_ada <= 975; v_din <= to_hexchar(dout[7:4]); end
976: begin v_ada <= 976; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h76 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
977: begin v_ada <= 977; v_din <= to_hexchar(dout[7:4]); end
978: begin v_ada <= 978; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h77 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
979: begin v_ada <= 979; v_din <= to_hexchar(dout[7:4]); end
980: begin v_ada <= 980; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h78 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
983: begin v_ada <= 983; v_din <= to_hexchar(dout[7:4]); end
984: begin v_ada <= 984; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h79 & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
985: begin v_ada <= 985; v_din <= to_hexchar(dout[7:4]); end
986: begin v_ada <= 986; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h7A & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
987: begin v_ada <= 987; v_din <= to_hexchar(dout[7:4]); end
988: begin v_ada <= 988; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h7B & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
989: begin v_ada <= 989; v_din <= to_hexchar(dout[7:4]); end
990: begin v_ada <= 990; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h7C & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
992: begin v_ada <= 992; v_din <= to_hexchar(dout[7:4]); end
993: begin v_ada <= 993; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h7D & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
994: begin v_ada <= 994; v_din <= to_hexchar(dout[7:4]); end
995: begin v_ada <= 995; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h7E & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
996: begin v_ada <= 996; v_din <= to_hexchar(dout[7:4]); end
997: begin v_ada <= 997; v_din <= to_hexchar(dout[3:0]);  adb <= operands[15:0] + 8'h7F & RAMW; state <= FETCH_REQ; fetch_stage <= FETCH_DATA; next_state <= SHOW_INFO_Z07; end
998: begin v_ada <= 998; v_din <= to_hexchar(dout[7:4]); end
999: begin v_ada <= 999; v_din <= to_hexchar(dout[3:0]); end
